`timescale 1ns / 10ps

module character_rom (
    input logic clk,
    input logic [9:0] char_addr,
    output logic [6:0] char_data_out
);
    logic [6:0] rom [0:1023];

    initial begin
        rom[0] = 7'h1C;
        rom[1] = 7'h22;
        rom[2] = 7'h2A;
        rom[3] = 7'h3A;
        rom[4] = 7'h1A;
        rom[5] = 7'h02;
        rom[6] = 7'h3C;
        rom[7] = 7'h00;
        rom[8] = 7'h08;
        rom[9] = 7'h14;
        rom[10] = 7'h22;
        rom[11] = 7'h22;
        rom[12] = 7'h3E;
        rom[13] = 7'h22;
        rom[14] = 7'h22;
        rom[15] = 7'h00;
        rom[16] = 7'h1E;
        rom[17] = 7'h22;
        rom[18] = 7'h22;
        rom[19] = 7'h1E;
        rom[20] = 7'h22;
        rom[21] = 7'h22;
        rom[22] = 7'h1E;
        rom[23] = 7'h00;
        rom[24] = 7'h1C;
        rom[25] = 7'h22;
        rom[26] = 7'h02;
        rom[27] = 7'h02;
        rom[28] = 7'h02;
        rom[29] = 7'h22;
        rom[30] = 7'h1C;
        rom[31] = 7'h00;
        rom[32] = 7'h1E;
        rom[33] = 7'h22;
        rom[34] = 7'h22;
        rom[35] = 7'h22;
        rom[36] = 7'h22;
        rom[37] = 7'h22;
        rom[38] = 7'h1E;
        rom[39] = 7'h00;
        rom[40] = 7'h3E;
        rom[41] = 7'h02;
        rom[42] = 7'h02;
        rom[43] = 7'h1E;
        rom[44] = 7'h02;
        rom[45] = 7'h02;
        rom[46] = 7'h3E;
        rom[47] = 7'h00;
        rom[48] = 7'h3E;
        rom[49] = 7'h02;
        rom[50] = 7'h02;
        rom[51] = 7'h1E;
        rom[52] = 7'h02;
        rom[53] = 7'h02;
        rom[54] = 7'h02;
        rom[55] = 7'h00;
        rom[56] = 7'h3C;
        rom[57] = 7'h02;
        rom[58] = 7'h02;
        rom[59] = 7'h02;
        rom[60] = 7'h32;
        rom[61] = 7'h22;
        rom[62] = 7'h3C;
        rom[63] = 7'h00;
        rom[64] = 7'h22;
        rom[65] = 7'h22;
        rom[66] = 7'h22;
        rom[67] = 7'h3E;
        rom[68] = 7'h22;
        rom[69] = 7'h22;
        rom[70] = 7'h22;
        rom[71] = 7'h00;
        rom[72] = 7'h1C;
        rom[73] = 7'h08;
        rom[74] = 7'h08;
        rom[75] = 7'h08;
        rom[76] = 7'h08;
        rom[77] = 7'h08;
        rom[78] = 7'h1C;
        rom[79] = 7'h00;
        rom[80] = 7'h20;
        rom[81] = 7'h20;
        rom[82] = 7'h20;
        rom[83] = 7'h20;
        rom[84] = 7'h20;
        rom[85] = 7'h22;
        rom[86] = 7'h1C;
        rom[87] = 7'h00;
        rom[88] = 7'h22;
        rom[89] = 7'h12;
        rom[90] = 7'h0A;
        rom[91] = 7'h06;
        rom[92] = 7'h0A;
        rom[93] = 7'h12;
        rom[94] = 7'h22;
        rom[95] = 7'h00;
        rom[96] = 7'h02;
        rom[97] = 7'h02;
        rom[98] = 7'h02;
        rom[99] = 7'h02;
        rom[100] = 7'h02;
        rom[101] = 7'h02;
        rom[102] = 7'h3E;
        rom[103] = 7'h00;
        rom[104] = 7'h22;
        rom[105] = 7'h36;
        rom[106] = 7'h2A;
        rom[107] = 7'h2A;
        rom[108] = 7'h22;
        rom[109] = 7'h22;
        rom[110] = 7'h22;
        rom[111] = 7'h00;
        rom[112] = 7'h22;
        rom[113] = 7'h22;
        rom[114] = 7'h26;
        rom[115] = 7'h2A;
        rom[116] = 7'h32;
        rom[117] = 7'h22;
        rom[118] = 7'h22;
        rom[119] = 7'h00;
        rom[120] = 7'h1C;
        rom[121] = 7'h22;
        rom[122] = 7'h22;
        rom[123] = 7'h22;
        rom[124] = 7'h22;
        rom[125] = 7'h22;
        rom[126] = 7'h1C;
        rom[127] = 7'h00;
        rom[128] = 7'h1E;
        rom[129] = 7'h22;
        rom[130] = 7'h22;
        rom[131] = 7'h1E;
        rom[132] = 7'h02;
        rom[133] = 7'h02;
        rom[134] = 7'h02;
        rom[135] = 7'h00;
        rom[136] = 7'h1C;
        rom[137] = 7'h22;
        rom[138] = 7'h22;
        rom[139] = 7'h22;
        rom[140] = 7'h2A;
        rom[141] = 7'h12;
        rom[142] = 7'h2C;
        rom[143] = 7'h00;
        rom[144] = 7'h1E;
        rom[145] = 7'h22;
        rom[146] = 7'h22;
        rom[147] = 7'h1E;
        rom[148] = 7'h0A;
        rom[149] = 7'h12;
        rom[150] = 7'h22;
        rom[151] = 7'h00;
        rom[152] = 7'h1C;
        rom[153] = 7'h22;
        rom[154] = 7'h02;
        rom[155] = 7'h1C;
        rom[156] = 7'h20;
        rom[157] = 7'h22;
        rom[158] = 7'h1C;
        rom[159] = 7'h00;
        rom[160] = 7'h3E;
        rom[161] = 7'h08;
        rom[162] = 7'h08;
        rom[163] = 7'h08;
        rom[164] = 7'h08;
        rom[165] = 7'h08;
        rom[166] = 7'h08;
        rom[167] = 7'h00;
        rom[168] = 7'h22;
        rom[169] = 7'h22;
        rom[170] = 7'h22;
        rom[171] = 7'h22;
        rom[172] = 7'h22;
        rom[173] = 7'h22;
        rom[174] = 7'h1C;
        rom[175] = 7'h00;
        rom[176] = 7'h22;
        rom[177] = 7'h22;
        rom[178] = 7'h22;
        rom[179] = 7'h22;
        rom[180] = 7'h22;
        rom[181] = 7'h14;
        rom[182] = 7'h08;
        rom[183] = 7'h00;
        rom[184] = 7'h22;
        rom[185] = 7'h22;
        rom[186] = 7'h22;
        rom[187] = 7'h2A;
        rom[188] = 7'h2A;
        rom[189] = 7'h36;
        rom[190] = 7'h22;
        rom[191] = 7'h00;
        rom[192] = 7'h22;
        rom[193] = 7'h22;
        rom[194] = 7'h14;
        rom[195] = 7'h08;
        rom[196] = 7'h14;
        rom[197] = 7'h22;
        rom[198] = 7'h22;
        rom[199] = 7'h00;
        rom[200] = 7'h22;
        rom[201] = 7'h22;
        rom[202] = 7'h14;
        rom[203] = 7'h08;
        rom[204] = 7'h08;
        rom[205] = 7'h08;
        rom[206] = 7'h08;
        rom[207] = 7'h00;
        rom[208] = 7'h3E;
        rom[209] = 7'h20;
        rom[210] = 7'h10;
        rom[211] = 7'h08;
        rom[212] = 7'h04;
        rom[213] = 7'h02;
        rom[214] = 7'h3E;
        rom[215] = 7'h00;
        rom[216] = 7'h3E;
        rom[217] = 7'h06;
        rom[218] = 7'h06;
        rom[219] = 7'h06;
        rom[220] = 7'h06;
        rom[221] = 7'h06;
        rom[222] = 7'h3E;
        rom[223] = 7'h00;
        rom[224] = 7'h00;
        rom[225] = 7'h02;
        rom[226] = 7'h04;
        rom[227] = 7'h08;
        rom[228] = 7'h10;
        rom[229] = 7'h20;
        rom[230] = 7'h00;
        rom[231] = 7'h00;
        rom[232] = 7'h3E;
        rom[233] = 7'h30;
        rom[234] = 7'h30;
        rom[235] = 7'h30;
        rom[236] = 7'h30;
        rom[237] = 7'h30;
        rom[238] = 7'h3E;
        rom[239] = 7'h00;
        rom[240] = 7'h00;
        rom[241] = 7'h00;
        rom[242] = 7'h08;
        rom[243] = 7'h14;
        rom[244] = 7'h22;
        rom[245] = 7'h00;
        rom[246] = 7'h00;
        rom[247] = 7'h00;
        rom[248] = 7'h00;
        rom[249] = 7'h00;
        rom[250] = 7'h00;
        rom[251] = 7'h00;
        rom[252] = 7'h00;
        rom[253] = 7'h00;
        rom[254] = 7'h00;
        rom[255] = 7'h7F;
        rom[256] = 7'h00;
        rom[257] = 7'h00;
        rom[258] = 7'h00;
        rom[259] = 7'h00;
        rom[260] = 7'h00;
        rom[261] = 7'h00;
        rom[262] = 7'h00;
        rom[263] = 7'h00;
        rom[264] = 7'h08;
        rom[265] = 7'h08;
        rom[266] = 7'h08;
        rom[267] = 7'h08;
        rom[268] = 7'h08;
        rom[269] = 7'h00;
        rom[270] = 7'h08;
        rom[271] = 7'h00;
        rom[272] = 7'h14;
        rom[273] = 7'h14;
        rom[274] = 7'h14;
        rom[275] = 7'h00;
        rom[276] = 7'h00;
        rom[277] = 7'h00;
        rom[278] = 7'h00;
        rom[279] = 7'h00;
        rom[280] = 7'h14;
        rom[281] = 7'h14;
        rom[282] = 7'h3E;
        rom[283] = 7'h14;
        rom[284] = 7'h3E;
        rom[285] = 7'h14;
        rom[286] = 7'h14;
        rom[287] = 7'h00;
        rom[288] = 7'h08;
        rom[289] = 7'h3C;
        rom[290] = 7'h0A;
        rom[291] = 7'h1C;
        rom[292] = 7'h28;
        rom[293] = 7'h1E;
        rom[294] = 7'h08;
        rom[295] = 7'h00;
        rom[296] = 7'h06;
        rom[297] = 7'h26;
        rom[298] = 7'h10;
        rom[299] = 7'h08;
        rom[300] = 7'h04;
        rom[301] = 7'h32;
        rom[302] = 7'h30;
        rom[303] = 7'h00;
        rom[304] = 7'h04;
        rom[305] = 7'h0A;
        rom[306] = 7'h0A;
        rom[307] = 7'h04;
        rom[308] = 7'h2A;
        rom[309] = 7'h12;
        rom[310] = 7'h2C;
        rom[311] = 7'h00;
        rom[312] = 7'h08;
        rom[313] = 7'h08;
        rom[314] = 7'h08;
        rom[315] = 7'h00;
        rom[316] = 7'h00;
        rom[317] = 7'h00;
        rom[318] = 7'h00;
        rom[319] = 7'h00;
        rom[320] = 7'h08;
        rom[321] = 7'h04;
        rom[322] = 7'h02;
        rom[323] = 7'h02;
        rom[324] = 7'h02;
        rom[325] = 7'h04;
        rom[326] = 7'h08;
        rom[327] = 7'h00;
        rom[328] = 7'h08;
        rom[329] = 7'h10;
        rom[330] = 7'h20;
        rom[331] = 7'h20;
        rom[332] = 7'h20;
        rom[333] = 7'h10;
        rom[334] = 7'h08;
        rom[335] = 7'h00;
        rom[336] = 7'h08;
        rom[337] = 7'h2A;
        rom[338] = 7'h1C;
        rom[339] = 7'h08;
        rom[340] = 7'h1C;
        rom[341] = 7'h2A;
        rom[342] = 7'h08;
        rom[343] = 7'h00;
        rom[344] = 7'h00;
        rom[345] = 7'h08;
        rom[346] = 7'h08;
        rom[347] = 7'h3E;
        rom[348] = 7'h08;
        rom[349] = 7'h08;
        rom[350] = 7'h00;
        rom[351] = 7'h00;
        rom[352] = 7'h00;
        rom[353] = 7'h00;
        rom[354] = 7'h00;
        rom[355] = 7'h00;
        rom[356] = 7'h08;
        rom[357] = 7'h08;
        rom[358] = 7'h04;
        rom[359] = 7'h00;
        rom[360] = 7'h00;
        rom[361] = 7'h00;
        rom[362] = 7'h00;
        rom[363] = 7'h3E;
        rom[364] = 7'h00;
        rom[365] = 7'h00;
        rom[366] = 7'h00;
        rom[367] = 7'h00;
        rom[368] = 7'h00;
        rom[369] = 7'h00;
        rom[370] = 7'h00;
        rom[371] = 7'h00;
        rom[372] = 7'h00;
        rom[373] = 7'h00;
        rom[374] = 7'h08;
        rom[375] = 7'h00;
        rom[376] = 7'h00;
        rom[377] = 7'h20;
        rom[378] = 7'h10;
        rom[379] = 7'h08;
        rom[380] = 7'h04;
        rom[381] = 7'h02;
        rom[382] = 7'h00;
        rom[383] = 7'h00;
        rom[384] = 7'h1C;
        rom[385] = 7'h22;
        rom[386] = 7'h32;
        rom[387] = 7'h2A;
        rom[388] = 7'h26;
        rom[389] = 7'h22;
        rom[390] = 7'h1C;
        rom[391] = 7'h00;
        rom[392] = 7'h08;
        rom[393] = 7'h0C;
        rom[394] = 7'h08;
        rom[395] = 7'h08;
        rom[396] = 7'h08;
        rom[397] = 7'h08;
        rom[398] = 7'h1C;
        rom[399] = 7'h00;
        rom[400] = 7'h1C;
        rom[401] = 7'h22;
        rom[402] = 7'h20;
        rom[403] = 7'h18;
        rom[404] = 7'h04;
        rom[405] = 7'h02;
        rom[406] = 7'h3E;
        rom[407] = 7'h00;
        rom[408] = 7'h3E;
        rom[409] = 7'h20;
        rom[410] = 7'h10;
        rom[411] = 7'h18;
        rom[412] = 7'h20;
        rom[413] = 7'h22;
        rom[414] = 7'h1C;
        rom[415] = 7'h00;
        rom[416] = 7'h10;
        rom[417] = 7'h18;
        rom[418] = 7'h14;
        rom[419] = 7'h12;
        rom[420] = 7'h3E;
        rom[421] = 7'h10;
        rom[422] = 7'h10;
        rom[423] = 7'h00;
        rom[424] = 7'h3E;
        rom[425] = 7'h02;
        rom[426] = 7'h1E;
        rom[427] = 7'h20;
        rom[428] = 7'h20;
        rom[429] = 7'h22;
        rom[430] = 7'h1C;
        rom[431] = 7'h00;
        rom[432] = 7'h38;
        rom[433] = 7'h04;
        rom[434] = 7'h02;
        rom[435] = 7'h1E;
        rom[436] = 7'h22;
        rom[437] = 7'h22;
        rom[438] = 7'h1C;
        rom[439] = 7'h00;
        rom[440] = 7'h3E;
        rom[441] = 7'h20;
        rom[442] = 7'h10;
        rom[443] = 7'h08;
        rom[444] = 7'h04;
        rom[445] = 7'h04;
        rom[446] = 7'h04;
        rom[447] = 7'h00;
        rom[448] = 7'h1C;
        rom[449] = 7'h22;
        rom[450] = 7'h22;
        rom[451] = 7'h1C;
        rom[452] = 7'h22;
        rom[453] = 7'h22;
        rom[454] = 7'h1C;
        rom[455] = 7'h00;
        rom[456] = 7'h1C;
        rom[457] = 7'h22;
        rom[458] = 7'h22;
        rom[459] = 7'h3C;
        rom[460] = 7'h20;
        rom[461] = 7'h10;
        rom[462] = 7'h0E;
        rom[463] = 7'h00;
        rom[464] = 7'h00;
        rom[465] = 7'h00;
        rom[466] = 7'h08;
        rom[467] = 7'h00;
        rom[468] = 7'h08;
        rom[469] = 7'h00;
        rom[470] = 7'h00;
        rom[471] = 7'h00;
        rom[472] = 7'h00;
        rom[473] = 7'h00;
        rom[474] = 7'h08;
        rom[475] = 7'h00;
        rom[476] = 7'h08;
        rom[477] = 7'h08;
        rom[478] = 7'h04;
        rom[479] = 7'h00;
        rom[480] = 7'h10;
        rom[481] = 7'h08;
        rom[482] = 7'h04;
        rom[483] = 7'h02;
        rom[484] = 7'h04;
        rom[485] = 7'h08;
        rom[486] = 7'h10;
        rom[487] = 7'h00;
        rom[488] = 7'h00;
        rom[489] = 7'h00;
        rom[490] = 7'h3E;
        rom[491] = 7'h00;
        rom[492] = 7'h3E;
        rom[493] = 7'h00;
        rom[494] = 7'h00;
        rom[495] = 7'h00;
        rom[496] = 7'h04;
        rom[497] = 7'h08;
        rom[498] = 7'h10;
        rom[499] = 7'h20;
        rom[500] = 7'h10;
        rom[501] = 7'h08;
        rom[502] = 7'h04;
        rom[503] = 7'h00;
        rom[504] = 7'h1C;
        rom[505] = 7'h22;
        rom[506] = 7'h10;
        rom[507] = 7'h08;
        rom[508] = 7'h08;
        rom[509] = 7'h00;
        rom[510] = 7'h08;
        rom[511] = 7'h00;
        rom[512] = 7'h1C;
        rom[513] = 7'h22;
        rom[514] = 7'h2A;
        rom[515] = 7'h3A;
        rom[516] = 7'h1A;
        rom[517] = 7'h02;
        rom[518] = 7'h3C;
        rom[519] = 7'h00;
        rom[520] = 7'h08;
        rom[521] = 7'h14;
        rom[522] = 7'h22;
        rom[523] = 7'h22;
        rom[524] = 7'h3E;
        rom[525] = 7'h22;
        rom[526] = 7'h22;
        rom[527] = 7'h00;
        rom[528] = 7'h1E;
        rom[529] = 7'h22;
        rom[530] = 7'h22;
        rom[531] = 7'h1E;
        rom[532] = 7'h22;
        rom[533] = 7'h22;
        rom[534] = 7'h1E;
        rom[535] = 7'h00;
        rom[536] = 7'h1C;
        rom[537] = 7'h22;
        rom[538] = 7'h02;
        rom[539] = 7'h02;
        rom[540] = 7'h02;
        rom[541] = 7'h22;
        rom[542] = 7'h1C;
        rom[543] = 7'h00;
        rom[544] = 7'h1E;
        rom[545] = 7'h22;
        rom[546] = 7'h22;
        rom[547] = 7'h22;
        rom[548] = 7'h22;
        rom[549] = 7'h22;
        rom[550] = 7'h1E;
        rom[551] = 7'h00;
        rom[552] = 7'h3E;
        rom[553] = 7'h02;
        rom[554] = 7'h02;
        rom[555] = 7'h1E;
        rom[556] = 7'h02;
        rom[557] = 7'h02;
        rom[558] = 7'h3E;
        rom[559] = 7'h00;
        rom[560] = 7'h3E;
        rom[561] = 7'h02;
        rom[562] = 7'h02;
        rom[563] = 7'h1E;
        rom[564] = 7'h02;
        rom[565] = 7'h02;
        rom[566] = 7'h02;
        rom[567] = 7'h00;
        rom[568] = 7'h3C;
        rom[569] = 7'h02;
        rom[570] = 7'h02;
        rom[571] = 7'h02;
        rom[572] = 7'h32;
        rom[573] = 7'h22;
        rom[574] = 7'h3C;
        rom[575] = 7'h00;
        rom[576] = 7'h22;
        rom[577] = 7'h22;
        rom[578] = 7'h22;
        rom[579] = 7'h3E;
        rom[580] = 7'h22;
        rom[581] = 7'h22;
        rom[582] = 7'h22;
        rom[583] = 7'h00;
        rom[584] = 7'h1C;
        rom[585] = 7'h08;
        rom[586] = 7'h08;
        rom[587] = 7'h08;
        rom[588] = 7'h08;
        rom[589] = 7'h08;
        rom[590] = 7'h1C;
        rom[591] = 7'h00;
        rom[592] = 7'h20;
        rom[593] = 7'h20;
        rom[594] = 7'h20;
        rom[595] = 7'h20;
        rom[596] = 7'h20;
        rom[597] = 7'h22;
        rom[598] = 7'h1C;
        rom[599] = 7'h00;
        rom[600] = 7'h22;
        rom[601] = 7'h12;
        rom[602] = 7'h0A;
        rom[603] = 7'h06;
        rom[604] = 7'h0A;
        rom[605] = 7'h12;
        rom[606] = 7'h22;
        rom[607] = 7'h00;
        rom[608] = 7'h02;
        rom[609] = 7'h02;
        rom[610] = 7'h02;
        rom[611] = 7'h02;
        rom[612] = 7'h02;
        rom[613] = 7'h02;
        rom[614] = 7'h3E;
        rom[615] = 7'h00;
        rom[616] = 7'h22;
        rom[617] = 7'h36;
        rom[618] = 7'h2A;
        rom[619] = 7'h2A;
        rom[620] = 7'h22;
        rom[621] = 7'h22;
        rom[622] = 7'h22;
        rom[623] = 7'h00;
        rom[624] = 7'h22;
        rom[625] = 7'h22;
        rom[626] = 7'h26;
        rom[627] = 7'h2A;
        rom[628] = 7'h32;
        rom[629] = 7'h22;
        rom[630] = 7'h22;
        rom[631] = 7'h00;
        rom[632] = 7'h1C;
        rom[633] = 7'h22;
        rom[634] = 7'h22;
        rom[635] = 7'h22;
        rom[636] = 7'h22;
        rom[637] = 7'h22;
        rom[638] = 7'h1C;
        rom[639] = 7'h00;
        rom[640] = 7'h1E;
        rom[641] = 7'h22;
        rom[642] = 7'h22;
        rom[643] = 7'h1E;
        rom[644] = 7'h02;
        rom[645] = 7'h02;
        rom[646] = 7'h02;
        rom[647] = 7'h00;
        rom[648] = 7'h1C;
        rom[649] = 7'h22;
        rom[650] = 7'h22;
        rom[651] = 7'h22;
        rom[652] = 7'h2A;
        rom[653] = 7'h12;
        rom[654] = 7'h2C;
        rom[655] = 7'h00;
        rom[656] = 7'h1E;
        rom[657] = 7'h22;
        rom[658] = 7'h22;
        rom[659] = 7'h1E;
        rom[660] = 7'h0A;
        rom[661] = 7'h12;
        rom[662] = 7'h22;
        rom[663] = 7'h00;
        rom[664] = 7'h1C;
        rom[665] = 7'h22;
        rom[666] = 7'h02;
        rom[667] = 7'h1C;
        rom[668] = 7'h20;
        rom[669] = 7'h22;
        rom[670] = 7'h1C;
        rom[671] = 7'h00;
        rom[672] = 7'h3E;
        rom[673] = 7'h08;
        rom[674] = 7'h08;
        rom[675] = 7'h08;
        rom[676] = 7'h08;
        rom[677] = 7'h08;
        rom[678] = 7'h08;
        rom[679] = 7'h00;
        rom[680] = 7'h22;
        rom[681] = 7'h22;
        rom[682] = 7'h22;
        rom[683] = 7'h22;
        rom[684] = 7'h22;
        rom[685] = 7'h22;
        rom[686] = 7'h1C;
        rom[687] = 7'h00;
        rom[688] = 7'h22;
        rom[689] = 7'h22;
        rom[690] = 7'h22;
        rom[691] = 7'h22;
        rom[692] = 7'h22;
        rom[693] = 7'h14;
        rom[694] = 7'h08;
        rom[695] = 7'h00;
        rom[696] = 7'h22;
        rom[697] = 7'h22;
        rom[698] = 7'h22;
        rom[699] = 7'h2A;
        rom[700] = 7'h2A;
        rom[701] = 7'h36;
        rom[702] = 7'h22;
        rom[703] = 7'h00;
        rom[704] = 7'h22;
        rom[705] = 7'h22;
        rom[706] = 7'h14;
        rom[707] = 7'h08;
        rom[708] = 7'h14;
        rom[709] = 7'h22;
        rom[710] = 7'h22;
        rom[711] = 7'h00;
        rom[712] = 7'h22;
        rom[713] = 7'h22;
        rom[714] = 7'h14;
        rom[715] = 7'h08;
        rom[716] = 7'h08;
        rom[717] = 7'h08;
        rom[718] = 7'h08;
        rom[719] = 7'h00;
        rom[720] = 7'h3E;
        rom[721] = 7'h20;
        rom[722] = 7'h10;
        rom[723] = 7'h08;
        rom[724] = 7'h04;
        rom[725] = 7'h02;
        rom[726] = 7'h3E;
        rom[727] = 7'h00;
        rom[728] = 7'h3E;
        rom[729] = 7'h06;
        rom[730] = 7'h06;
        rom[731] = 7'h06;
        rom[732] = 7'h06;
        rom[733] = 7'h06;
        rom[734] = 7'h3E;
        rom[735] = 7'h00;
        rom[736] = 7'h00;
        rom[737] = 7'h02;
        rom[738] = 7'h04;
        rom[739] = 7'h08;
        rom[740] = 7'h10;
        rom[741] = 7'h20;
        rom[742] = 7'h00;
        rom[743] = 7'h00;
        rom[744] = 7'h3E;
        rom[745] = 7'h30;
        rom[746] = 7'h30;
        rom[747] = 7'h30;
        rom[748] = 7'h30;
        rom[749] = 7'h30;
        rom[750] = 7'h3E;
        rom[751] = 7'h00;
        rom[752] = 7'h00;
        rom[753] = 7'h00;
        rom[754] = 7'h08;
        rom[755] = 7'h14;
        rom[756] = 7'h22;
        rom[757] = 7'h00;
        rom[758] = 7'h00;
        rom[759] = 7'h00;
        rom[760] = 7'h00;
        rom[761] = 7'h00;
        rom[762] = 7'h00;
        rom[763] = 7'h00;
        rom[764] = 7'h00;
        rom[765] = 7'h00;
        rom[766] = 7'h00;
        rom[767] = 7'h7F;
        rom[768] = 7'h04;
        rom[769] = 7'h08;
        rom[770] = 7'h10;
        rom[771] = 7'h00;
        rom[772] = 7'h00;
        rom[773] = 7'h00;
        rom[774] = 7'h00;
        rom[775] = 7'h00;
        rom[776] = 7'h00;
        rom[777] = 7'h00;
        rom[778] = 7'h1C;
        rom[779] = 7'h20;
        rom[780] = 7'h3C;
        rom[781] = 7'h22;
        rom[782] = 7'h3C;
        rom[783] = 7'h00;
        rom[784] = 7'h02;
        rom[785] = 7'h02;
        rom[786] = 7'h1E;
        rom[787] = 7'h22;
        rom[788] = 7'h22;
        rom[789] = 7'h22;
        rom[790] = 7'h1E;
        rom[791] = 7'h00;
        rom[792] = 7'h00;
        rom[793] = 7'h00;
        rom[794] = 7'h3C;
        rom[795] = 7'h02;
        rom[796] = 7'h02;
        rom[797] = 7'h02;
        rom[798] = 7'h3C;
        rom[799] = 7'h00;
        rom[800] = 7'h20;
        rom[801] = 7'h20;
        rom[802] = 7'h3C;
        rom[803] = 7'h22;
        rom[804] = 7'h22;
        rom[805] = 7'h22;
        rom[806] = 7'h3C;
        rom[807] = 7'h00;
        rom[808] = 7'h00;
        rom[809] = 7'h00;
        rom[810] = 7'h1C;
        rom[811] = 7'h22;
        rom[812] = 7'h3E;
        rom[813] = 7'h02;
        rom[814] = 7'h3C;
        rom[815] = 7'h00;
        rom[816] = 7'h18;
        rom[817] = 7'h24;
        rom[818] = 7'h04;
        rom[819] = 7'h1E;
        rom[820] = 7'h04;
        rom[821] = 7'h04;
        rom[822] = 7'h04;
        rom[823] = 7'h00;
        rom[824] = 7'h00;
        rom[825] = 7'h00;
        rom[826] = 7'h1C;
        rom[827] = 7'h22;
        rom[828] = 7'h22;
        rom[829] = 7'h3C;
        rom[830] = 7'h20;
        rom[831] = 7'h1C;
        rom[832] = 7'h02;
        rom[833] = 7'h02;
        rom[834] = 7'h1E;
        rom[835] = 7'h22;
        rom[836] = 7'h22;
        rom[837] = 7'h22;
        rom[838] = 7'h22;
        rom[839] = 7'h00;
        rom[840] = 7'h08;
        rom[841] = 7'h00;
        rom[842] = 7'h0C;
        rom[843] = 7'h08;
        rom[844] = 7'h08;
        rom[845] = 7'h08;
        rom[846] = 7'h1C;
        rom[847] = 7'h00;
        rom[848] = 7'h10;
        rom[849] = 7'h00;
        rom[850] = 7'h18;
        rom[851] = 7'h10;
        rom[852] = 7'h10;
        rom[853] = 7'h10;
        rom[854] = 7'h12;
        rom[855] = 7'h0C;
        rom[856] = 7'h02;
        rom[857] = 7'h02;
        rom[858] = 7'h22;
        rom[859] = 7'h12;
        rom[860] = 7'h0E;
        rom[861] = 7'h12;
        rom[862] = 7'h22;
        rom[863] = 7'h00;
        rom[864] = 7'h0C;
        rom[865] = 7'h08;
        rom[866] = 7'h08;
        rom[867] = 7'h08;
        rom[868] = 7'h08;
        rom[869] = 7'h08;
        rom[870] = 7'h1C;
        rom[871] = 7'h00;
        rom[872] = 7'h00;
        rom[873] = 7'h00;
        rom[874] = 7'h36;
        rom[875] = 7'h2A;
        rom[876] = 7'h2A;
        rom[877] = 7'h2A;
        rom[878] = 7'h22;
        rom[879] = 7'h00;
        rom[880] = 7'h00;
        rom[881] = 7'h00;
        rom[882] = 7'h1E;
        rom[883] = 7'h22;
        rom[884] = 7'h22;
        rom[885] = 7'h22;
        rom[886] = 7'h22;
        rom[887] = 7'h00;
        rom[888] = 7'h00;
        rom[889] = 7'h00;
        rom[890] = 7'h1C;
        rom[891] = 7'h22;
        rom[892] = 7'h22;
        rom[893] = 7'h22;
        rom[894] = 7'h1C;
        rom[895] = 7'h00;
        rom[896] = 7'h00;
        rom[897] = 7'h00;
        rom[898] = 7'h1E;
        rom[899] = 7'h22;
        rom[900] = 7'h22;
        rom[901] = 7'h1E;
        rom[902] = 7'h02;
        rom[903] = 7'h02;
        rom[904] = 7'h00;
        rom[905] = 7'h00;
        rom[906] = 7'h3C;
        rom[907] = 7'h22;
        rom[908] = 7'h22;
        rom[909] = 7'h3C;
        rom[910] = 7'h20;
        rom[911] = 7'h20;
        rom[912] = 7'h00;
        rom[913] = 7'h00;
        rom[914] = 7'h3A;
        rom[915] = 7'h06;
        rom[916] = 7'h02;
        rom[917] = 7'h02;
        rom[918] = 7'h02;
        rom[919] = 7'h00;
        rom[920] = 7'h00;
        rom[921] = 7'h00;
        rom[922] = 7'h3C;
        rom[923] = 7'h02;
        rom[924] = 7'h1C;
        rom[925] = 7'h20;
        rom[926] = 7'h1E;
        rom[927] = 7'h00;
        rom[928] = 7'h04;
        rom[929] = 7'h04;
        rom[930] = 7'h1E;
        rom[931] = 7'h04;
        rom[932] = 7'h04;
        rom[933] = 7'h24;
        rom[934] = 7'h18;
        rom[935] = 7'h00;
        rom[936] = 7'h00;
        rom[937] = 7'h00;
        rom[938] = 7'h22;
        rom[939] = 7'h22;
        rom[940] = 7'h22;
        rom[941] = 7'h32;
        rom[942] = 7'h2C;
        rom[943] = 7'h00;
        rom[944] = 7'h00;
        rom[945] = 7'h00;
        rom[946] = 7'h22;
        rom[947] = 7'h22;
        rom[948] = 7'h22;
        rom[949] = 7'h14;
        rom[950] = 7'h08;
        rom[951] = 7'h00;
        rom[952] = 7'h00;
        rom[953] = 7'h00;
        rom[954] = 7'h22;
        rom[955] = 7'h22;
        rom[956] = 7'h2A;
        rom[957] = 7'h2A;
        rom[958] = 7'h36;
        rom[959] = 7'h00;
        rom[960] = 7'h00;
        rom[961] = 7'h00;
        rom[962] = 7'h22;
        rom[963] = 7'h14;
        rom[964] = 7'h08;
        rom[965] = 7'h14;
        rom[966] = 7'h22;
        rom[967] = 7'h00;
        rom[968] = 7'h00;
        rom[969] = 7'h00;
        rom[970] = 7'h22;
        rom[971] = 7'h22;
        rom[972] = 7'h22;
        rom[973] = 7'h3C;
        rom[974] = 7'h20;
        rom[975] = 7'h1C;
        rom[976] = 7'h00;
        rom[977] = 7'h00;
        rom[978] = 7'h3E;
        rom[979] = 7'h10;
        rom[980] = 7'h08;
        rom[981] = 7'h04;
        rom[982] = 7'h3E;
        rom[983] = 7'h00;
        rom[984] = 7'h38;
        rom[985] = 7'h0C;
        rom[986] = 7'h0C;
        rom[987] = 7'h06;
        rom[988] = 7'h0C;
        rom[989] = 7'h0C;
        rom[990] = 7'h38;
        rom[991] = 7'h00;
        rom[992] = 7'h08;
        rom[993] = 7'h08;
        rom[994] = 7'h08;
        rom[995] = 7'h08;
        rom[996] = 7'h08;
        rom[997] = 7'h08;
        rom[998] = 7'h08;
        rom[999] = 7'h08;
        rom[1000] = 7'h0E;
        rom[1001] = 7'h18;
        rom[1002] = 7'h18;
        rom[1003] = 7'h30;
        rom[1004] = 7'h18;
        rom[1005] = 7'h18;
        rom[1006] = 7'h0E;
        rom[1007] = 7'h00;
        rom[1008] = 7'h2C;
        rom[1009] = 7'h1A;
        rom[1010] = 7'h00;
        rom[1011] = 7'h00;
        rom[1012] = 7'h00;
        rom[1013] = 7'h00;
        rom[1014] = 7'h00;
        rom[1015] = 7'h00;
        rom[1016] = 7'h00;
        rom[1017] = 7'h2A;
        rom[1018] = 7'h14;
        rom[1019] = 7'h2A;
        rom[1020] = 7'h14;
        rom[1021] = 7'h2A;
        rom[1022] = 7'h00;
        rom[1023] = 7'h00;
    end

    always_ff @(posedge clk) begin
        char_data_out <= rom[char_addr];        
    end

endmodule