module apple2_ram #(
    parameter ADDR_WIDTH = 16,
    parameter DATA_WIDTH = 8
)(
    // CLOCK SIGNALS we need
    input logic CPUCLK, VGACLK,

    // KEYBOARD
    input logic [7:0] decoded,
    input logic oflag,
    // ADDRESS PORTS
    input logic [ADDR_WIDTH - 1:0] CPUADDR, VGAADDR,
    
    // ENABLE PORTs for CPU WRITE
    input logic CPU_WEN, 
    
    // DATA INPUTS
    input logic [7:0] DSTORE,

    // DATA OUTPUTS
    output logic [7:0] CPU_DOUT, VGA_DOUT
);

(* ram_style = "block" *) reg [DATA_WIDTH-1:0] mem [0:(1 << ADDR_WIDTH) - 1];

// CPU Port (write/read)
always_ff @(posedge CPUCLK) begin
    if(CPU_WEN) begin
         mem[CPUADDR] <= DSTORE; 
    end else begin
        CPU_DOUT <= mem[CPUADDR];
    end
end

// VGA Port (read-only)
always_ff @(posedge VGACLK) begin
    VGA_DOUT <= mem[VGAADDR];
end

initial begin
    for(integer i = 16'h0000; i < 16'hD000; i++) begin
      mem[i] = 8'b0;
    end
    mem[16'h0000] = 8'h00;
mem[16'h0001] = 8'h9C;
mem[16'h0002] = 8'h00;
mem[16'h0003] = 8'h08;
mem[16'h0004] = 8'h3A;
mem[16'h0005] = 8'h03;
mem[16'h0006] = 8'h00;
mem[16'h0007] = 8'h00;
mem[16'h0008] = 8'h00;
mem[16'h0009] = 8'hC0;
mem[16'h000A] = 8'h60;
mem[16'h000B] = 8'h01;
mem[16'h000C] = 8'h05;
mem[16'h000D] = 8'h00;
mem[16'h000E] = 8'h00;
mem[16'h000F] = 8'h6B;
mem[16'h0010] = 8'h00;
mem[16'h0011] = 8'h9C;
mem[16'h0012] = 8'h00;
mem[16'h0013] = 8'h04;
mem[16'h0014] = 8'h00;
mem[16'h0015] = 8'h00;
mem[16'h0016] = 8'h00;
mem[16'h0017] = 8'h00;
mem[16'h0018] = 8'hFF;
mem[16'h0019] = 8'h0C;
mem[16'h001A] = 8'h00;
mem[16'h001B] = 8'h56;
mem[16'h001C] = 8'hFF;
mem[16'h001D] = 8'hFF;
mem[16'h001E] = 8'h00;
mem[16'h001F] = 8'h00;
mem[16'h0020] = 8'h00;
mem[16'h0021] = 8'h28;
mem[16'h0022] = 8'h00;
mem[16'h0023] = 8'h18;
mem[16'h0024] = 8'h26;
mem[16'h0025] = 8'h17;
mem[16'h0026] = 8'h70;
mem[16'h0027] = 8'h06;
mem[16'h0028] = 8'h80;
mem[16'h0029] = 8'h04;
mem[16'h002A] = 8'hF5;
mem[16'h002B] = 8'h43;
mem[16'h002C] = 8'h00;
mem[16'h002D] = 8'h00;
mem[16'h002E] = 8'hE8;
mem[16'h002F] = 8'h01;
mem[16'h0030] = 8'hFE;
mem[16'h0031] = 8'h00;
mem[16'h0032] = 8'hFF;
mem[16'h0033] = 8'hAA;
mem[16'h0034] = 8'h05;
mem[16'h0035] = 8'h28;
mem[16'h0036] = 8'h09;
mem[16'h0037] = 8'h03;
mem[16'h0038] = 8'h1B;
mem[16'h0039] = 8'hFD;
mem[16'h003A] = 8'hFF;
mem[16'h003B] = 8'hBF;
mem[16'h003C] = 8'h00;
mem[16'h003D] = 8'h9C;
mem[16'h003E] = 8'h00;
mem[16'h003F] = 8'h9C;
mem[16'h0040] = 8'h00;
mem[16'h0041] = 8'h9C;
mem[16'h0042] = 8'hA2;
mem[16'h0043] = 8'h5B;
mem[16'h0044] = 8'h82;
mem[16'h0045] = 8'h98;
mem[16'h0046] = 8'h62;
mem[16'h0047] = 8'hD8;
mem[16'h0048] = 8'h00;
mem[16'h0049] = 8'hB7;
mem[16'h004A] = 8'h00;
mem[16'h004B] = 8'h00;
mem[16'h004C] = 8'hFF;
mem[16'h004D] = 8'hFF;
mem[16'h004E] = 8'h14;
mem[16'h004F] = 8'h07;
mem[16'h0050] = 8'h26;
mem[16'h0051] = 8'hFF;
mem[16'h0052] = 8'h41;
mem[16'h0053] = 8'h02;
mem[16'h0054] = 8'h00;
mem[16'h0055] = 8'h00;
mem[16'h0056] = 8'hBC;
mem[16'h0057] = 8'h7E;
mem[16'h0058] = 8'hFF;
mem[16'h0059] = 8'hD0;
mem[16'h005A] = 8'h2F;
mem[16'h005B] = 8'h00;
mem[16'h005C] = 8'h00;
mem[16'h005D] = 8'hFF;
mem[16'h005E] = 8'hD1;
mem[16'h005F] = 8'h4D;
mem[16'h0060] = 8'hA5;
mem[16'h0061] = 8'h00;
mem[16'h0062] = 8'h19;
mem[16'h0063] = 8'h00;
mem[16'h0064] = 8'h00;
mem[16'h0065] = 8'h00;
mem[16'h0066] = 8'h0E;
mem[16'h0067] = 8'h38;
mem[16'h0068] = 8'h00;
mem[16'h0069] = 8'h00;
mem[16'h006A] = 8'h00;
mem[16'h006B] = 8'h00;
mem[16'h006C] = 8'h00;
mem[16'h006D] = 8'h00;
mem[16'h006E] = 8'h01;
mem[16'h006F] = 8'h33;
mem[16'h0070] = 8'h08;
mem[16'h0071] = 8'hFF;
mem[16'h0072] = 8'h00;
mem[16'h0073] = 8'h05;
mem[16'h0074] = 8'h60;
mem[16'h0075] = 8'h18;
mem[16'h0076] = 8'h27;
mem[16'h0077] = 8'h01;
mem[16'h0078] = 8'h7F;
mem[16'h0079] = 8'h41;
mem[16'h007A] = 8'h83;
mem[16'h007B] = 8'h7E;
mem[16'h007C] = 8'h83;
mem[16'h007D] = 8'hC1;
mem[16'h007E] = 8'hDA;
mem[16'h007F] = 8'h88;
mem[16'h0080] = 8'h95;
mem[16'h0081] = 8'hFF;
mem[16'h0082] = 8'h00;
mem[16'h0083] = 8'h00;
mem[16'h0084] = 8'hFF;
mem[16'h0085] = 8'h00;
mem[16'h0086] = 8'h00;
mem[16'h0087] = 8'h00;
mem[16'h0088] = 8'h00;
mem[16'h0089] = 8'h00;
mem[16'h008A] = 8'h00;
mem[16'h008B] = 8'h00;
mem[16'h008C] = 8'hFF;
mem[16'h008D] = 8'hFF;
mem[16'h008E] = 8'h00;
mem[16'h008F] = 8'h03;
mem[16'h0090] = 8'h4C;
mem[16'h0091] = 8'h64;
mem[16'h0092] = 8'h00;
mem[16'h0093] = 8'h00;
mem[16'h0094] = 8'hFF;
mem[16'h0095] = 8'hFF;
mem[16'h0096] = 8'h00;
mem[16'h0097] = 8'h00;
mem[16'h0098] = 8'hFF;
mem[16'h0099] = 8'h00;
mem[16'h009A] = 8'h00;
mem[16'h009B] = 8'h00;
mem[16'h009C] = 8'h00;
mem[16'h009D] = 8'h88;
mem[16'h009E] = 8'hFF;
mem[16'h009F] = 8'hFF;
mem[16'h00A0] = 8'hFF;
mem[16'h00A1] = 8'h69;
mem[16'h00A2] = 8'hFF;
mem[16'h00A3] = 8'h00;
mem[16'h00A4] = 8'h00;
mem[16'h00A5] = 8'hD0;
mem[16'h00A6] = 8'hD1;
mem[16'h00A7] = 8'hFF;
mem[16'h00A8] = 8'hFF;
mem[16'h00A9] = 8'h69;
mem[16'h00AA] = 8'hFF;
mem[16'h00AB] = 8'hFF;
mem[16'h00AC] = 8'h00;
mem[16'h00AD] = 8'h09;
mem[16'h00AE] = 8'h08;
mem[16'h00AF] = 8'h04;
mem[16'h00B0] = 8'h08;
mem[16'h00B1] = 8'hE6;
mem[16'h00B2] = 8'hB8;
mem[16'h00B3] = 8'hD0;
mem[16'h00B4] = 8'h02;
mem[16'h00B5] = 8'hE6;
mem[16'h00B6] = 8'hB9;
mem[16'h00B7] = 8'hAD;
mem[16'h00B8] = 8'h05;
mem[16'h00B9] = 8'h02;
mem[16'h00BA] = 8'hC9;
mem[16'h00BB] = 8'h3A;
mem[16'h00BC] = 8'hB0;
mem[16'h00BD] = 8'h0A;
mem[16'h00BE] = 8'hC9;
mem[16'h00BF] = 8'h20;
mem[16'h00C0] = 8'hF0;
mem[16'h00C1] = 8'hEF;
mem[16'h00C2] = 8'h38;
mem[16'h00C3] = 8'hE9;
mem[16'h00C4] = 8'h30;
mem[16'h00C5] = 8'h38;
mem[16'h00C6] = 8'hE9;
mem[16'h00C7] = 8'hD0;
mem[16'h00C8] = 8'h60;
mem[16'h00C9] = 8'h80;
mem[16'h00CA] = 8'h4F;
mem[16'h00CB] = 8'hC7;
mem[16'h00CC] = 8'h52;
mem[16'h00CD] = 8'hFF;
mem[16'h00CE] = 8'h00;
mem[16'h00CF] = 8'h00;
mem[16'h00D0] = 8'hFF;
mem[16'h00D1] = 8'hFF;
mem[16'h00D2] = 8'h00;
mem[16'h00D3] = 8'h00;
mem[16'h00D4] = 8'hFF;
mem[16'h00D5] = 8'hFF;
mem[16'h00D6] = 8'h00;
mem[16'h00D7] = 8'h00;
mem[16'h00D8] = 8'h00;
mem[16'h00D9] = 8'hFF;
mem[16'h00DA] = 8'h00;
mem[16'h00DB] = 8'h00;
mem[16'h00DC] = 8'hFF;
mem[16'h00DD] = 8'hFF;
mem[16'h00DE] = 8'h00;
mem[16'h00DF] = 8'h00;
mem[16'h00E0] = 8'hFF;
mem[16'h00E1] = 8'hFF;
mem[16'h00E2] = 8'h00;
mem[16'h00E3] = 8'h00;
mem[16'h00E4] = 8'hFF;
mem[16'h00E5] = 8'hFF;
mem[16'h00E6] = 8'h00;
mem[16'h00E7] = 8'h00;
mem[16'h00E8] = 8'hFF;
mem[16'h00E9] = 8'hFF;
mem[16'h00EA] = 8'h00;
mem[16'h00EB] = 8'h00;
mem[16'h00EC] = 8'hFF;
mem[16'h00ED] = 8'hFF;
mem[16'h00EE] = 8'h00;
mem[16'h00EF] = 8'h00;
mem[16'h00F0] = 8'hFF;
mem[16'h00F1] = 8'h01;
mem[16'h00F2] = 8'h00;
mem[16'h00F3] = 8'h00;
mem[16'h00F4] = 8'hFF;
mem[16'h00F5] = 8'hFF;
mem[16'h00F6] = 8'h00;
mem[16'h00F7] = 8'h00;
mem[16'h00F8] = 8'hF8;
mem[16'h00F9] = 8'hFF;
mem[16'h00FA] = 8'h00;
mem[16'h00FB] = 8'h00;
mem[16'h00FC] = 8'hFF;
mem[16'h00FD] = 8'hFF;
mem[16'h00FE] = 8'h00;
mem[16'h00FF] = 8'h10;
mem[16'h0100] = 8'h00;
mem[16'h0101] = 8'hFF;
mem[16'h0102] = 8'h00;
mem[16'h0103] = 8'h00;
mem[16'h0104] = 8'h00;
mem[16'h0105] = 8'hFF;
mem[16'h0106] = 8'h00;
mem[16'h0107] = 8'h00;
mem[16'h0108] = 8'h00;
mem[16'h0109] = 8'hFF;
mem[16'h010A] = 8'h00;
mem[16'h010B] = 8'h00;
mem[16'h010C] = 8'h00;
mem[16'h010D] = 8'hFF;
mem[16'h010E] = 8'h00;
mem[16'h010F] = 8'h00;
mem[16'h0110] = 8'h00;
mem[16'h0111] = 8'hFF;
mem[16'h0112] = 8'h00;
mem[16'h0113] = 8'h00;
mem[16'h0114] = 8'h00;
mem[16'h0115] = 8'hFF;
mem[16'h0116] = 8'h00;
mem[16'h0117] = 8'h00;
mem[16'h0118] = 8'h00;
mem[16'h0119] = 8'hFF;
mem[16'h011A] = 8'h00;
mem[16'h011B] = 8'h00;
mem[16'h011C] = 8'h00;
mem[16'h011D] = 8'hFF;
mem[16'h011E] = 8'h00;
mem[16'h011F] = 8'h00;
mem[16'h0120] = 8'h00;
mem[16'h0121] = 8'hFF;
mem[16'h0122] = 8'h00;
mem[16'h0123] = 8'h00;
mem[16'h0124] = 8'h00;
mem[16'h0125] = 8'hFF;
mem[16'h0126] = 8'h00;
mem[16'h0127] = 8'h00;
mem[16'h0128] = 8'h00;
mem[16'h0129] = 8'hFF;
mem[16'h012A] = 8'h00;
mem[16'h012B] = 8'h00;
mem[16'h012C] = 8'h00;
mem[16'h012D] = 8'hFF;
mem[16'h012E] = 8'h00;
mem[16'h012F] = 8'h00;
mem[16'h0130] = 8'h00;
mem[16'h0131] = 8'hFF;
mem[16'h0132] = 8'h00;
mem[16'h0133] = 8'h00;
mem[16'h0134] = 8'h00;
mem[16'h0135] = 8'hFF;
mem[16'h0136] = 8'h00;
mem[16'h0137] = 8'h00;
mem[16'h0138] = 8'h00;
mem[16'h0139] = 8'hFF;
mem[16'h013A] = 8'h00;
mem[16'h013B] = 8'h00;
mem[16'h013C] = 8'h00;
mem[16'h013D] = 8'hFF;
mem[16'h013E] = 8'h00;
mem[16'h013F] = 8'h00;
mem[16'h0140] = 8'h00;
mem[16'h0141] = 8'hFF;
mem[16'h0142] = 8'h00;
mem[16'h0143] = 8'h00;
mem[16'h0144] = 8'h00;
mem[16'h0145] = 8'hFF;
mem[16'h0146] = 8'h00;
mem[16'h0147] = 8'h00;
mem[16'h0148] = 8'h00;
mem[16'h0149] = 8'hFF;
mem[16'h014A] = 8'h00;
mem[16'h014B] = 8'h00;
mem[16'h014C] = 8'h00;
mem[16'h014D] = 8'hFF;
mem[16'h014E] = 8'h00;
mem[16'h014F] = 8'h00;
mem[16'h0150] = 8'h00;
mem[16'h0151] = 8'hFF;
mem[16'h0152] = 8'h00;
mem[16'h0153] = 8'h00;
mem[16'h0154] = 8'h00;
mem[16'h0155] = 8'hFF;
mem[16'h0156] = 8'h00;
mem[16'h0157] = 8'h00;
mem[16'h0158] = 8'h00;
mem[16'h0159] = 8'hFF;
mem[16'h015A] = 8'h00;
mem[16'h015B] = 8'h00;
mem[16'h015C] = 8'h00;
mem[16'h015D] = 8'hFF;
mem[16'h015E] = 8'h00;
mem[16'h015F] = 8'h00;
mem[16'h0160] = 8'h00;
mem[16'h0161] = 8'hFF;
mem[16'h0162] = 8'h00;
mem[16'h0163] = 8'h00;
mem[16'h0164] = 8'h00;
mem[16'h0165] = 8'hFF;
mem[16'h0166] = 8'h00;
mem[16'h0167] = 8'h00;
mem[16'h0168] = 8'h00;
mem[16'h0169] = 8'hFF;
mem[16'h016A] = 8'h00;
mem[16'h016B] = 8'h00;
mem[16'h016C] = 8'h00;
mem[16'h016D] = 8'hFF;
mem[16'h016E] = 8'h00;
mem[16'h016F] = 8'h00;
mem[16'h0170] = 8'h00;
mem[16'h0171] = 8'hFF;
mem[16'h0172] = 8'h00;
mem[16'h0173] = 8'h00;
mem[16'h0174] = 8'h00;
mem[16'h0175] = 8'hFF;
mem[16'h0176] = 8'h00;
mem[16'h0177] = 8'h00;
mem[16'h0178] = 8'h00;
mem[16'h0179] = 8'hFF;
mem[16'h017A] = 8'h00;
mem[16'h017B] = 8'h00;
mem[16'h017C] = 8'h00;
mem[16'h017D] = 8'hFF;
mem[16'h017E] = 8'h00;
mem[16'h017F] = 8'h00;
mem[16'h0180] = 8'h00;
mem[16'h0181] = 8'hFF;
mem[16'h0182] = 8'h00;
mem[16'h0183] = 8'h00;
mem[16'h0184] = 8'h00;
mem[16'h0185] = 8'hFF;
mem[16'h0186] = 8'h00;
mem[16'h0187] = 8'h00;
mem[16'h0188] = 8'h00;
mem[16'h0189] = 8'hFF;
mem[16'h018A] = 8'h00;
mem[16'h018B] = 8'h00;
mem[16'h018C] = 8'h00;
mem[16'h018D] = 8'hFF;
mem[16'h018E] = 8'h00;
mem[16'h018F] = 8'h00;
mem[16'h0190] = 8'h00;
mem[16'h0191] = 8'hFF;
mem[16'h0192] = 8'h00;
mem[16'h0193] = 8'h00;
mem[16'h0194] = 8'h00;
mem[16'h0195] = 8'hFF;
mem[16'h0196] = 8'h00;
mem[16'h0197] = 8'h00;
mem[16'h0198] = 8'h00;
mem[16'h0199] = 8'hFF;
mem[16'h019A] = 8'h00;
mem[16'h019B] = 8'h00;
mem[16'h019C] = 8'h00;
mem[16'h019D] = 8'hFF;
mem[16'h019E] = 8'h00;
mem[16'h019F] = 8'h00;
mem[16'h01A0] = 8'h00;
mem[16'h01A1] = 8'hFF;
mem[16'h01A2] = 8'h00;
mem[16'h01A3] = 8'h00;
mem[16'h01A4] = 8'h00;
mem[16'h01A5] = 8'hFF;
mem[16'h01A6] = 8'h00;
mem[16'h01A7] = 8'h00;
mem[16'h01A8] = 8'h00;
mem[16'h01A9] = 8'hFF;
mem[16'h01AA] = 8'h00;
mem[16'h01AB] = 8'h00;
mem[16'h01AC] = 8'h00;
mem[16'h01AD] = 8'hFF;
mem[16'h01AE] = 8'h00;
mem[16'h01AF] = 8'h00;
mem[16'h01B0] = 8'h00;
mem[16'h01B1] = 8'hFF;
mem[16'h01B2] = 8'h00;
mem[16'h01B3] = 8'h00;
mem[16'h01B4] = 8'h00;
mem[16'h01B5] = 8'hFF;
mem[16'h01B6] = 8'h00;
mem[16'h01B7] = 8'h00;
mem[16'h01B8] = 8'h00;
mem[16'h01B9] = 8'hFF;
mem[16'h01BA] = 8'h00;
mem[16'h01BB] = 8'h00;
mem[16'h01BC] = 8'h00;
mem[16'h01BD] = 8'hFF;
mem[16'h01BE] = 8'h00;
mem[16'h01BF] = 8'h00;
mem[16'h01C0] = 8'h00;
mem[16'h01C1] = 8'hFF;
mem[16'h01C2] = 8'h00;
mem[16'h01C3] = 8'h00;
mem[16'h01C4] = 8'h00;
mem[16'h01C5] = 8'hFF;
mem[16'h01C6] = 8'h00;
mem[16'h01C7] = 8'h00;
mem[16'h01C8] = 8'h00;
mem[16'h01C9] = 8'hFF;
mem[16'h01CA] = 8'h39;
mem[16'h01CB] = 8'hB5;
mem[16'h01CC] = 8'h38;
mem[16'h01CD] = 8'hB7;
mem[16'h01CE] = 8'hDA;
mem[16'h01CF] = 8'hB6;
mem[16'h01D0] = 8'h4F;
mem[16'h01D1] = 8'hB6;
mem[16'h01D2] = 8'h5F;
mem[16'h01D3] = 8'hBF;
mem[16'h01D4] = 8'h20;
mem[16'h01D5] = 8'hB4;
mem[16'h01D6] = 8'h09;
mem[16'h01D7] = 8'h00;
mem[16'h01D8] = 8'hB0;
mem[16'h01D9] = 8'h02;
mem[16'h01DA] = 8'h10;
mem[16'h01DB] = 8'hCF;
mem[16'h01DC] = 8'h5F;
mem[16'h01DD] = 8'h0B;
mem[16'h01DE] = 8'h40;
mem[16'h01DF] = 8'h84;
mem[16'h01E0] = 8'hFF;
mem[16'h01E1] = 8'h26;
mem[16'h01E2] = 8'hFC;
mem[16'h01E3] = 8'hA0;
mem[16'h01E4] = 8'h37;
mem[16'h01E5] = 8'h6D;
mem[16'h01E6] = 8'h00;
mem[16'h01E7] = 8'h36;
mem[16'h01E8] = 8'h83;
mem[16'h01E9] = 8'hBA;
mem[16'h01EA] = 8'h82;
mem[16'h01EB] = 8'hDA;
mem[16'h01EC] = 8'h6F;
mem[16'h01ED] = 8'h55;
mem[16'h01EE] = 8'h40;
mem[16'h01EF] = 8'hCF;
mem[16'h01F0] = 8'h5F;
mem[16'h01F1] = 8'h0B;
mem[16'h01F2] = 8'h40;
mem[16'h01F3] = 8'h69;
mem[16'h01F4] = 8'h00;
mem[16'h01F5] = 8'h6F;
mem[16'h01F6] = 8'h00;
mem[16'h01F7] = 8'h22;
mem[16'h01F8] = 8'h00;
mem[16'h01F9] = 8'hC1;
mem[16'h01FA] = 8'h00;
mem[16'h01FB] = 8'h00;
mem[16'h01FC] = 8'h00;
mem[16'h01FD] = 8'h01;
mem[16'h01FE] = 8'h00;
mem[16'h01FF] = 8'h37;
mem[16'h0200] = 8'hB9;
mem[16'h0201] = 8'hC3;
mem[16'h0202] = 8'hB0;
mem[16'h0203] = 8'hB0;
mem[16'h0204] = 8'hC7;
mem[16'h0205] = 8'h8D;
mem[16'h0206] = 8'hC6;
mem[16'h0207] = 8'hB5;
mem[16'h0208] = 8'hB9;
mem[16'h0209] = 8'h8D;
mem[16'h020A] = 8'hD8;
mem[16'h020B] = 8'h8D;
mem[16'h020C] = 8'h8D;
mem[16'h020D] = 8'hB1;
mem[16'h020E] = 8'h8D;
mem[16'h020F] = 8'hAC;
mem[16'h0210] = 8'h00;
mem[16'h0211] = 8'hA4;
mem[16'h0212] = 8'h00;
mem[16'h0213] = 8'hB0;
mem[16'h0214] = 8'h00;
mem[16'h0215] = 8'hB0;
mem[16'h0216] = 8'h00;
mem[16'h0217] = 8'hCC;
mem[16'h0218] = 8'h00;
mem[16'h0219] = 8'hB2;
mem[16'h021A] = 8'h00;
mem[16'h021B] = 8'hB0;
mem[16'h021C] = 8'h00;
mem[16'h021D] = 8'h8D;
mem[16'h021E] = 8'h00;
mem[16'h021F] = 8'h00;
mem[16'h0220] = 8'h00;
mem[16'h0221] = 8'hFF;
mem[16'h0222] = 8'h00;
mem[16'h0223] = 8'h02;
mem[16'h0224] = 8'h00;
mem[16'h0225] = 8'hFF;
mem[16'h0226] = 8'h00;
mem[16'h0227] = 8'h02;
mem[16'h0228] = 8'h00;
mem[16'h0229] = 8'hFF;
mem[16'h022A] = 8'h00;
mem[16'h022B] = 8'h02;
mem[16'h022C] = 8'h00;
mem[16'h022D] = 8'hFF;
mem[16'h022E] = 8'h00;
mem[16'h022F] = 8'h02;
mem[16'h0230] = 8'h00;
mem[16'h0231] = 8'hFF;
mem[16'h0232] = 8'h00;
mem[16'h0233] = 8'h00;
mem[16'h0234] = 8'h00;
mem[16'h0235] = 8'hFF;
mem[16'h0236] = 8'h00;
mem[16'h0237] = 8'h00;
mem[16'h0238] = 8'h00;
mem[16'h0239] = 8'hFF;
mem[16'h023A] = 8'h00;
mem[16'h023B] = 8'h00;
mem[16'h023C] = 8'h00;
mem[16'h023D] = 8'hFF;
mem[16'h023E] = 8'h00;
mem[16'h023F] = 8'h00;
mem[16'h0240] = 8'h00;
mem[16'h0241] = 8'hFF;
mem[16'h0242] = 8'h00;
mem[16'h0243] = 8'h00;
mem[16'h0244] = 8'h00;
mem[16'h0245] = 8'hFF;
mem[16'h0246] = 8'h00;
mem[16'h0247] = 8'h00;
mem[16'h0248] = 8'h00;
mem[16'h0249] = 8'hFF;
mem[16'h024A] = 8'h00;
mem[16'h024B] = 8'h00;
mem[16'h024C] = 8'h00;
mem[16'h024D] = 8'hFF;
mem[16'h024E] = 8'h00;
mem[16'h024F] = 8'h00;
mem[16'h0250] = 8'h00;
mem[16'h0251] = 8'hFF;
mem[16'h0252] = 8'h00;
mem[16'h0253] = 8'h00;
mem[16'h0254] = 8'h00;
mem[16'h0255] = 8'hFF;
mem[16'h0256] = 8'h00;
mem[16'h0257] = 8'h00;
mem[16'h0258] = 8'h00;
mem[16'h0259] = 8'hFF;
mem[16'h025A] = 8'h00;
mem[16'h025B] = 8'h00;
mem[16'h025C] = 8'h00;
mem[16'h025D] = 8'hFF;
mem[16'h025E] = 8'h00;
mem[16'h025F] = 8'h00;
mem[16'h0260] = 8'h00;
mem[16'h0261] = 8'hFF;
mem[16'h0262] = 8'h00;
mem[16'h0263] = 8'h00;
mem[16'h0264] = 8'h00;
mem[16'h0265] = 8'hFF;
mem[16'h0266] = 8'h00;
mem[16'h0267] = 8'h00;
mem[16'h0268] = 8'h00;
mem[16'h0269] = 8'hFF;
mem[16'h026A] = 8'h00;
mem[16'h026B] = 8'h00;
mem[16'h026C] = 8'h00;
mem[16'h026D] = 8'hFF;
mem[16'h026E] = 8'h00;
mem[16'h026F] = 8'h00;
mem[16'h0270] = 8'h00;
mem[16'h0271] = 8'hFF;
mem[16'h0272] = 8'h00;
mem[16'h0273] = 8'h00;
mem[16'h0274] = 8'h00;
mem[16'h0275] = 8'hFF;
mem[16'h0276] = 8'h00;
mem[16'h0277] = 8'h00;
mem[16'h0278] = 8'h00;
mem[16'h0279] = 8'hFF;
mem[16'h027A] = 8'h00;
mem[16'h027B] = 8'h00;
mem[16'h027C] = 8'h00;
mem[16'h027D] = 8'hFF;
mem[16'h027E] = 8'h00;
mem[16'h027F] = 8'h00;
mem[16'h0280] = 8'h00;
mem[16'h0281] = 8'hFF;
mem[16'h0282] = 8'h00;
mem[16'h0283] = 8'h00;
mem[16'h0284] = 8'h00;
mem[16'h0285] = 8'hFF;
mem[16'h0286] = 8'h00;
mem[16'h0287] = 8'h00;
mem[16'h0288] = 8'h00;
mem[16'h0289] = 8'hFF;
mem[16'h028A] = 8'h00;
mem[16'h028B] = 8'h00;
mem[16'h028C] = 8'h00;
mem[16'h028D] = 8'hFF;
mem[16'h028E] = 8'h00;
mem[16'h028F] = 8'h02;
mem[16'h0290] = 8'h00;
mem[16'h0291] = 8'hFF;
mem[16'h0292] = 8'h00;
mem[16'h0293] = 8'h00;
mem[16'h0294] = 8'h00;
mem[16'h0295] = 8'hFF;
mem[16'h0296] = 8'h00;
mem[16'h0297] = 8'h00;
mem[16'h0298] = 8'h00;
mem[16'h0299] = 8'hFF;
mem[16'h029A] = 8'h00;
mem[16'h029B] = 8'h00;
mem[16'h029C] = 8'h00;
mem[16'h029D] = 8'hFF;
mem[16'h029E] = 8'h00;
mem[16'h029F] = 8'h00;
mem[16'h02A0] = 8'h00;
mem[16'h02A1] = 8'hFF;
mem[16'h02A2] = 8'h00;
mem[16'h02A3] = 8'h02;
mem[16'h02A4] = 8'h00;
mem[16'h02A5] = 8'hFF;
mem[16'h02A6] = 8'h00;
mem[16'h02A7] = 8'h02;
mem[16'h02A8] = 8'h00;
mem[16'h02A9] = 8'hFF;
mem[16'h02AA] = 8'h00;
mem[16'h02AB] = 8'h00;
mem[16'h02AC] = 8'h00;
mem[16'h02AD] = 8'hFF;
mem[16'h02AE] = 8'h00;
mem[16'h02AF] = 8'h02;
mem[16'h02B0] = 8'h00;
mem[16'h02B1] = 8'hFF;
mem[16'h02B2] = 8'h00;
mem[16'h02B3] = 8'h00;
mem[16'h02B4] = 8'h00;
mem[16'h02B5] = 8'hFF;
mem[16'h02B6] = 8'h00;
mem[16'h02B7] = 8'h00;
mem[16'h02B8] = 8'h00;
mem[16'h02B9] = 8'hFF;
mem[16'h02BA] = 8'h00;
mem[16'h02BB] = 8'h00;
mem[16'h02BC] = 8'h00;
mem[16'h02BD] = 8'hFF;
mem[16'h02BE] = 8'h00;
mem[16'h02BF] = 8'h00;
mem[16'h02C0] = 8'h00;
mem[16'h02C1] = 8'hFF;
mem[16'h02C2] = 8'h00;
mem[16'h02C3] = 8'h00;
mem[16'h02C4] = 8'h00;
mem[16'h02C5] = 8'hFF;
mem[16'h02C6] = 8'h00;
mem[16'h02C7] = 8'h00;
mem[16'h02C8] = 8'h00;
mem[16'h02C9] = 8'hFF;
mem[16'h02CA] = 8'h00;
mem[16'h02CB] = 8'h00;
mem[16'h02CC] = 8'h00;
mem[16'h02CD] = 8'hFF;
mem[16'h02CE] = 8'h00;
mem[16'h02CF] = 8'h00;
mem[16'h02D0] = 8'h00;
mem[16'h02D1] = 8'hFF;
mem[16'h02D2] = 8'h00;
mem[16'h02D3] = 8'h00;
mem[16'h02D4] = 8'h00;
mem[16'h02D5] = 8'hFF;
mem[16'h02D6] = 8'h00;
mem[16'h02D7] = 8'h00;
mem[16'h02D8] = 8'h00;
mem[16'h02D9] = 8'hFF;
mem[16'h02DA] = 8'h00;
mem[16'h02DB] = 8'h00;
mem[16'h02DC] = 8'h00;
mem[16'h02DD] = 8'hFF;
mem[16'h02DE] = 8'h00;
mem[16'h02DF] = 8'h00;
mem[16'h02E0] = 8'h00;
mem[16'h02E1] = 8'hFF;
mem[16'h02E2] = 8'h00;
mem[16'h02E3] = 8'h00;
mem[16'h02E4] = 8'h00;
mem[16'h02E5] = 8'hFF;
mem[16'h02E6] = 8'h00;
mem[16'h02E7] = 8'h00;
mem[16'h02E8] = 8'h00;
mem[16'h02E9] = 8'hFF;
mem[16'h02EA] = 8'h00;
mem[16'h02EB] = 8'h00;
mem[16'h02EC] = 8'h00;
mem[16'h02ED] = 8'hFF;
mem[16'h02EE] = 8'h00;
mem[16'h02EF] = 8'h00;
mem[16'h02F0] = 8'h00;
mem[16'h02F1] = 8'hFF;
mem[16'h02F2] = 8'h00;
mem[16'h02F3] = 8'h00;
mem[16'h02F4] = 8'h00;
mem[16'h02F5] = 8'hFF;
mem[16'h02F6] = 8'h00;
mem[16'h02F7] = 8'h00;
mem[16'h02F8] = 8'h00;
mem[16'h02F9] = 8'hFF;
mem[16'h02FA] = 8'h00;
mem[16'h02FB] = 8'h00;
mem[16'h02FC] = 8'h00;
mem[16'h02FD] = 8'hFF;
mem[16'h02FE] = 8'h00;
mem[16'h02FF] = 8'h00;
mem[16'h0300] = 8'hA0;
mem[16'h0301] = 8'h03;
mem[16'h0302] = 8'h84;
mem[16'h0303] = 8'h37;
mem[16'h0304] = 8'hA0;
mem[16'h0305] = 8'h09;
mem[16'h0306] = 8'h84;
mem[16'h0307] = 8'h36;
mem[16'h0308] = 8'h60;
mem[16'h0309] = 8'h48;
mem[16'h030A] = 8'h84;
mem[16'h030B] = 8'h4E;
mem[16'h030C] = 8'hC9;
mem[16'h030D] = 8'h8D;
mem[16'h030E] = 8'hF0;
mem[16'h030F] = 8'h68;
mem[16'h0310] = 8'hA5;
mem[16'h0311] = 8'h25;
mem[16'h0312] = 8'h4A;
mem[16'h0313] = 8'h29;
mem[16'h0314] = 8'h03;
mem[16'h0315] = 8'h09;
mem[16'h0316] = 8'h20;
mem[16'h0317] = 8'h85;
mem[16'h0318] = 8'h2B;
mem[16'h0319] = 8'hA5;
mem[16'h031A] = 8'h25;
mem[16'h031B] = 8'h6A;
mem[16'h031C] = 8'h08;
mem[16'h031D] = 8'h0A;
mem[16'h031E] = 8'h29;
mem[16'h031F] = 8'h18;
mem[16'h0320] = 8'h85;
mem[16'h0321] = 8'h2A;
mem[16'h0322] = 8'h0A;
mem[16'h0323] = 8'h0A;
mem[16'h0324] = 8'h05;
mem[16'h0325] = 8'h2A;
mem[16'h0326] = 8'h0A;
mem[16'h0327] = 8'h28;
mem[16'h0328] = 8'h6A;
mem[16'h0329] = 8'h18;
mem[16'h032A] = 8'h65;
mem[16'h032B] = 8'h24;
mem[16'h032C] = 8'h85;
mem[16'h032D] = 8'h2A;
mem[16'h032E] = 8'h68;
mem[16'h032F] = 8'h29;
mem[16'h0330] = 8'h7F;
mem[16'h0331] = 8'h48;
mem[16'h0332] = 8'hA9;
mem[16'h0333] = 8'h00;
mem[16'h0334] = 8'h85;
mem[16'h0335] = 8'h27;
mem[16'h0336] = 8'h68;
mem[16'h0337] = 8'h48;
mem[16'h0338] = 8'h2A;
mem[16'h0339] = 8'h26;
mem[16'h033A] = 8'h27;
mem[16'h033B] = 8'h2A;
mem[16'h033C] = 8'h26;
mem[16'h033D] = 8'h27;
mem[16'h033E] = 8'h2A;
mem[16'h033F] = 8'h26;
mem[16'h0340] = 8'h27;
mem[16'h0341] = 8'h85;
mem[16'h0342] = 8'h26;
mem[16'h0343] = 8'hA5;
mem[16'h0344] = 8'h27;
mem[16'h0345] = 8'h18;
mem[16'h0346] = 8'h69;
mem[16'h0347] = 8'h04;
mem[16'h0348] = 8'h85;
mem[16'h0349] = 8'h27;
mem[16'h034A] = 8'hA0;
mem[16'h034B] = 8'h00;
mem[16'h034C] = 8'hB1;
mem[16'h034D] = 8'h26;
mem[16'h034E] = 8'h48;
mem[16'h034F] = 8'h84;
mem[16'h0350] = 8'h4F;
mem[16'h0351] = 8'hA0;
mem[16'h0352] = 8'h00;
mem[16'h0353] = 8'h51;
mem[16'h0354] = 8'h2A;
mem[16'h0355] = 8'h91;
mem[16'h0356] = 8'h2A;
mem[16'h0357] = 8'hA5;
mem[16'h0358] = 8'h2B;
mem[16'h0359] = 8'hEA;
mem[16'h035A] = 8'hEA;
mem[16'h035B] = 8'h85;
mem[16'h035C] = 8'h2B;
mem[16'h035D] = 8'h68;
mem[16'h035E] = 8'h51;
mem[16'h035F] = 8'h2A;
mem[16'h0360] = 8'hEA;
mem[16'h0361] = 8'hEA;
mem[16'h0362] = 8'hA4;
mem[16'h0363] = 8'h4F;
mem[16'h0364] = 8'hA5;
mem[16'h0365] = 8'h2B;
mem[16'h0366] = 8'h18;
mem[16'h0367] = 8'h69;
mem[16'h0368] = 8'h04;
mem[16'h0369] = 8'h85;
mem[16'h036A] = 8'h2B;
mem[16'h036B] = 8'hC8;
mem[16'h036C] = 8'hC0;
mem[16'h036D] = 8'h08;
mem[16'h036E] = 8'hD0;
mem[16'h036F] = 8'hDC;
mem[16'h0370] = 8'hE6;
mem[16'h0371] = 8'h24;
mem[16'h0372] = 8'hA5;
mem[16'h0373] = 8'h24;
mem[16'h0374] = 8'hC5;
mem[16'h0375] = 8'h21;
mem[16'h0376] = 8'h90;
mem[16'h0377] = 8'h10;
mem[16'h0378] = 8'hA5;
mem[16'h0379] = 8'h20;
mem[16'h037A] = 8'h85;
mem[16'h037B] = 8'h24;
mem[16'h037C] = 8'hE6;
mem[16'h037D] = 8'h25;
mem[16'h037E] = 8'hA5;
mem[16'h037F] = 8'h25;
mem[16'h0380] = 8'hC5;
mem[16'h0381] = 8'h23;
mem[16'h0382] = 8'h90;
mem[16'h0383] = 8'h04;
mem[16'h0384] = 8'hA5;
mem[16'h0385] = 8'h22;
mem[16'h0386] = 8'h85;
mem[16'h0387] = 8'h25;
mem[16'h0388] = 8'hA4;
mem[16'h0389] = 8'h4E;
mem[16'h038A] = 8'h68;
mem[16'h038B] = 8'h60;
mem[16'h038C] = 8'hFF;
mem[16'h038D] = 8'hFF;
mem[16'h038E] = 8'h00;
mem[16'h038F] = 8'h00;
mem[16'h0390] = 8'hFF;
mem[16'h0391] = 8'hFF;
mem[16'h0392] = 8'h00;
mem[16'h0393] = 8'h00;
mem[16'h0394] = 8'hFF;
mem[16'h0395] = 8'hFF;
mem[16'h0396] = 8'h00;
mem[16'h0397] = 8'h00;
mem[16'h0398] = 8'hFF;
mem[16'h0399] = 8'hFF;
mem[16'h039A] = 8'h00;
mem[16'h039B] = 8'h00;
mem[16'h039C] = 8'hFF;
mem[16'h039D] = 8'hFF;
mem[16'h039E] = 8'h00;
mem[16'h039F] = 8'h00;
mem[16'h03A0] = 8'hFF;
mem[16'h03A1] = 8'hFF;
mem[16'h03A2] = 8'h00;
mem[16'h03A3] = 8'h00;
mem[16'h03A4] = 8'hFF;
mem[16'h03A5] = 8'hFF;
mem[16'h03A6] = 8'h00;
mem[16'h03A7] = 8'h00;
mem[16'h03A8] = 8'hFF;
mem[16'h03A9] = 8'hFF;
mem[16'h03AA] = 8'h00;
mem[16'h03AB] = 8'h00;
mem[16'h03AC] = 8'hFF;
mem[16'h03AD] = 8'hFF;
mem[16'h03AE] = 8'h00;
mem[16'h03AF] = 8'h00;
mem[16'h03B0] = 8'hFF;
mem[16'h03B1] = 8'hFF;
mem[16'h03B2] = 8'h00;
mem[16'h03B3] = 8'h00;
mem[16'h03B4] = 8'hFF;
mem[16'h03B5] = 8'hFF;
mem[16'h03B6] = 8'h00;
mem[16'h03B7] = 8'h00;
mem[16'h03B8] = 8'hFF;
mem[16'h03B9] = 8'hFF;
mem[16'h03BA] = 8'h00;
mem[16'h03BB] = 8'h00;
mem[16'h03BC] = 8'hFF;
mem[16'h03BD] = 8'hFF;
mem[16'h03BE] = 8'h00;
mem[16'h03BF] = 8'h00;
mem[16'h03C0] = 8'h00;
mem[16'h03C1] = 8'h00;
mem[16'h03C2] = 8'h00;
mem[16'h03C3] = 8'h00;
mem[16'h03C4] = 8'h00;
mem[16'h03C5] = 8'h00;
mem[16'h03C6] = 8'h00;
mem[16'h03C7] = 8'h00;
mem[16'h03C8] = 8'h00;
mem[16'h03C9] = 8'h00;
mem[16'h03CA] = 8'h00;
mem[16'h03CB] = 8'h00;
mem[16'h03CC] = 8'hB6;
mem[16'h03CD] = 8'h00;
mem[16'h03CE] = 8'h00;
mem[16'h03CF] = 8'h00;
mem[16'h03D0] = 8'h4C;
mem[16'h03D1] = 8'hBF;
mem[16'h03D2] = 8'h9D;
mem[16'h03D3] = 8'h4C;
mem[16'h03D4] = 8'h84;
mem[16'h03D5] = 8'h9D;
mem[16'h03D6] = 8'h4C;
mem[16'h03D7] = 8'hFD;
mem[16'h03D8] = 8'hAA;
mem[16'h03D9] = 8'h4C;
mem[16'h03DA] = 8'hB5;
mem[16'h03DB] = 8'hB7;
mem[16'h03DC] = 8'hAD;
mem[16'h03DD] = 8'h0F;
mem[16'h03DE] = 8'h9D;
mem[16'h03DF] = 8'hAC;
mem[16'h03E0] = 8'h0E;
mem[16'h03E1] = 8'h9D;
mem[16'h03E2] = 8'h60;
mem[16'h03E3] = 8'hAD;
mem[16'h03E4] = 8'hC2;
mem[16'h03E5] = 8'hAA;
mem[16'h03E6] = 8'hAC;
mem[16'h03E7] = 8'hC1;
mem[16'h03E8] = 8'hAA;
mem[16'h03E9] = 8'h60;
mem[16'h03EA] = 8'h4C;
mem[16'h03EB] = 8'h51;
mem[16'h03EC] = 8'hA8;
mem[16'h03ED] = 8'hEA;
mem[16'h03EE] = 8'hEA;
mem[16'h03EF] = 8'h4C;
mem[16'h03F0] = 8'h59;
mem[16'h03F1] = 8'hFA;
mem[16'h03F2] = 8'h43;
mem[16'h03F3] = 8'h00;
mem[16'h03F4] = 8'hAE;
mem[16'h03F5] = 8'h4C;
mem[16'h03F6] = 8'h58;
mem[16'h03F7] = 8'hFF;
mem[16'h03F8] = 8'h4C;
mem[16'h03F9] = 8'h65;
mem[16'h03FA] = 8'hFF;
mem[16'h03FB] = 8'h4C;
mem[16'h03FC] = 8'h65;
mem[16'h03FD] = 8'hFF;
mem[16'h03FE] = 8'h65;
mem[16'h03FF] = 8'hFF;
mem[16'h0400] = 8'h00;
mem[16'h0401] = 8'hFF;
mem[16'h0402] = 8'hFF;
mem[16'h0403] = 8'h00;
mem[16'h0404] = 8'h00;
mem[16'h0405] = 8'hFF;
mem[16'h0406] = 8'hFF;
mem[16'h0407] = 8'h00;
mem[16'h0408] = 8'h00;
mem[16'h0409] = 8'hFF;
mem[16'h040A] = 8'hFF;
mem[16'h040B] = 8'h00;
mem[16'h040C] = 8'h00;
mem[16'h040D] = 8'hFF;
mem[16'h040E] = 8'hFF;
mem[16'h040F] = 8'h00;
mem[16'h0410] = 8'h00;
mem[16'h0411] = 8'hFF;
mem[16'h0412] = 8'hFF;
mem[16'h0413] = 8'h00;
mem[16'h0414] = 8'h00;
mem[16'h0415] = 8'hFF;
mem[16'h0416] = 8'hFF;
mem[16'h0417] = 8'h00;
mem[16'h0418] = 8'h00;
mem[16'h0419] = 8'hFF;
mem[16'h041A] = 8'hFF;
mem[16'h041B] = 8'h00;
mem[16'h041C] = 8'h00;
mem[16'h041D] = 8'hFF;
mem[16'h041E] = 8'hFF;
mem[16'h041F] = 8'h00;
mem[16'h0420] = 8'h00;
mem[16'h0421] = 8'hFF;
mem[16'h0422] = 8'hFF;
mem[16'h0423] = 8'h00;
mem[16'h0424] = 8'h00;
mem[16'h0425] = 8'hFF;
mem[16'h0426] = 8'hFF;
mem[16'h0427] = 8'h00;
mem[16'h0428] = 8'h00;
mem[16'h0429] = 8'hFF;
mem[16'h042A] = 8'hFF;
mem[16'h042B] = 8'h00;
mem[16'h042C] = 8'h00;
mem[16'h042D] = 8'hFF;
mem[16'h042E] = 8'hFF;
mem[16'h042F] = 8'h00;
mem[16'h0430] = 8'h00;
mem[16'h0431] = 8'hFF;
mem[16'h0432] = 8'hFF;
mem[16'h0433] = 8'h00;
mem[16'h0434] = 8'h00;
mem[16'h0435] = 8'hFF;
mem[16'h0436] = 8'hFF;
mem[16'h0437] = 8'h00;
mem[16'h0438] = 8'h00;
mem[16'h0439] = 8'h14;
mem[16'h043A] = 8'h22;
mem[16'h043B] = 8'h22;
mem[16'h043C] = 8'h22;
mem[16'h043D] = 8'h41;
mem[16'h043E] = 8'h7F;
mem[16'h043F] = 8'h08;
mem[16'h0440] = 8'h10;
mem[16'h0441] = 8'h08;
mem[16'h0442] = 8'h04;
mem[16'h0443] = 8'h7E;
mem[16'h0444] = 8'h04;
mem[16'h0445] = 8'h08;
mem[16'h0446] = 8'h10;
mem[16'h0447] = 8'h00;
mem[16'h0448] = 8'h08;
mem[16'h0449] = 8'h10;
mem[16'h044A] = 8'h20;
mem[16'h044B] = 8'h7E;
mem[16'h044C] = 8'h20;
mem[16'h044D] = 8'h10;
mem[16'h044E] = 8'h08;
mem[16'h044F] = 8'h00;
mem[16'h0450] = 8'h08;
mem[16'h0451] = 8'h08;
mem[16'h0452] = 8'h08;
mem[16'h0453] = 8'h49;
mem[16'h0454] = 8'h2A;
mem[16'h0455] = 8'h1C;
mem[16'h0456] = 8'h08;
mem[16'h0457] = 8'h00;
mem[16'h0458] = 8'h08;
mem[16'h0459] = 8'h1C;
mem[16'h045A] = 8'h2A;
mem[16'h045B] = 8'h49;
mem[16'h045C] = 8'h08;
mem[16'h045D] = 8'h08;
mem[16'h045E] = 8'h08;
mem[16'h045F] = 8'h00;
mem[16'h0460] = 8'h08;
mem[16'h0461] = 8'h49;
mem[16'h0462] = 8'h2A;
mem[16'h0463] = 8'h1C;
mem[16'h0464] = 8'h49;
mem[16'h0465] = 8'h2A;
mem[16'h0466] = 8'h1C;
mem[16'h0467] = 8'h08;
mem[16'h0468] = 8'h40;
mem[16'h0469] = 8'h60;
mem[16'h046A] = 8'h70;
mem[16'h046B] = 8'h78;
mem[16'h046C] = 8'h70;
mem[16'h046D] = 8'h60;
mem[16'h046E] = 8'h40;
mem[16'h046F] = 8'h00;
mem[16'h0470] = 8'h40;
mem[16'h0471] = 8'h40;
mem[16'h0472] = 8'h20;
mem[16'h0473] = 8'h20;
mem[16'h0474] = 8'h13;
mem[16'h0475] = 8'h14;
mem[16'h0476] = 8'h0C;
mem[16'h0477] = 8'h08;
mem[16'h0478] = 8'h1A;
mem[16'h0479] = 8'h00;
mem[16'h047A] = 8'h00;
mem[16'h047B] = 8'h7C;
mem[16'h047C] = 8'h2A;
mem[16'h047D] = 8'h28;
mem[16'h047E] = 8'h34;
mem[16'h047F] = 8'h00;
mem[16'h0480] = 8'h36;
mem[16'h0481] = 8'h7F;
mem[16'h0482] = 8'h7F;
mem[16'h0483] = 8'h7F;
mem[16'h0484] = 8'h3E;
mem[16'h0485] = 8'h1C;
mem[16'h0486] = 8'h08;
mem[16'h0487] = 8'h00;
mem[16'h0488] = 8'h08;
mem[16'h0489] = 8'h1C;
mem[16'h048A] = 8'h3E;
mem[16'h048B] = 8'h7F;
mem[16'h048C] = 8'h3E;
mem[16'h048D] = 8'h1C;
mem[16'h048E] = 8'h08;
mem[16'h048F] = 8'h00;
mem[16'h0490] = 8'h08;
mem[16'h0491] = 8'h1C;
mem[16'h0492] = 8'h3E;
mem[16'h0493] = 8'h7F;
mem[16'h0494] = 8'h7F;
mem[16'h0495] = 8'h2A;
mem[16'h0496] = 8'h08;
mem[16'h0497] = 8'h00;
mem[16'h0498] = 8'h08;
mem[16'h0499] = 8'h1C;
mem[16'h049A] = 8'h1C;
mem[16'h049B] = 8'h2A;
mem[16'h049C] = 8'h7F;
mem[16'h049D] = 8'h7F;
mem[16'h049E] = 8'h2A;
mem[16'h049F] = 8'h08;
mem[16'h04A0] = 8'h3E;
mem[16'h04A1] = 8'h08;
mem[16'h04A2] = 8'h08;
mem[16'h04A3] = 8'h22;
mem[16'h04A4] = 8'h36;
mem[16'h04A5] = 8'h2A;
mem[16'h04A6] = 8'h22;
mem[16'h04A7] = 8'h00;
mem[16'h04A8] = 8'h00;
mem[16'h04A9] = 8'h22;
mem[16'h04AA] = 8'h14;
mem[16'h04AB] = 8'h08;
mem[16'h04AC] = 8'h14;
mem[16'h04AD] = 8'h22;
mem[16'h04AE] = 8'h00;
mem[16'h04AF] = 8'h00;
mem[16'h04B0] = 8'h04;
mem[16'h04B1] = 8'h0E;
mem[16'h04B2] = 8'h04;
mem[16'h04B3] = 8'h04;
mem[16'h04B4] = 8'h00;
mem[16'h04B5] = 8'h00;
mem[16'h04B6] = 8'h00;
mem[16'h04B7] = 8'h00;
mem[16'h04B8] = 8'h00;
mem[16'h04B9] = 8'h08;
mem[16'h04BA] = 8'h00;
mem[16'h04BB] = 8'h3E;
mem[16'h04BC] = 8'h00;
mem[16'h04BD] = 8'h08;
mem[16'h04BE] = 8'h00;
mem[16'h04BF] = 8'h00;
mem[16'h04C0] = 8'h18;
mem[16'h04C1] = 8'h24;
mem[16'h04C2] = 8'h08;
mem[16'h04C3] = 8'h14;
mem[16'h04C4] = 8'h08;
mem[16'h04C5] = 8'h12;
mem[16'h04C6] = 8'h0C;
mem[16'h04C7] = 8'h00;
mem[16'h04C8] = 8'h10;
mem[16'h04C9] = 8'h38;
mem[16'h04CA] = 8'h04;
mem[16'h04CB] = 8'h04;
mem[16'h04CC] = 8'h38;
mem[16'h04CD] = 8'h10;
mem[16'h04CE] = 8'h00;
mem[16'h04CF] = 8'h00;
mem[16'h04D0] = 8'h08;
mem[16'h04D1] = 8'h1C;
mem[16'h04D2] = 8'h08;
mem[16'h04D3] = 8'h1C;
mem[16'h04D4] = 8'h3E;
mem[16'h04D5] = 8'h1C;
mem[16'h04D6] = 8'h3E;
mem[16'h04D7] = 8'h7F;
mem[16'h04D8] = 8'h08;
mem[16'h04D9] = 8'h3E;
mem[16'h04DA] = 8'h1C;
mem[16'h04DB] = 8'h08;
mem[16'h04DC] = 8'h1C;
mem[16'h04DD] = 8'h1C;
mem[16'h04DE] = 8'h3E;
mem[16'h04DF] = 8'h7F;
mem[16'h04E0] = 8'h00;
mem[16'h04E1] = 8'h2A;
mem[16'h04E2] = 8'h3E;
mem[16'h04E3] = 8'h1C;
mem[16'h04E4] = 8'h1C;
mem[16'h04E5] = 8'h1C;
mem[16'h04E6] = 8'h3E;
mem[16'h04E7] = 8'h7F;
mem[16'h04E8] = 8'h00;
mem[16'h04E9] = 8'h10;
mem[16'h04EA] = 8'h3C;
mem[16'h04EB] = 8'h3E;
mem[16'h04EC] = 8'h18;
mem[16'h04ED] = 8'h0C;
mem[16'h04EE] = 8'h1E;
mem[16'h04EF] = 8'h3F;
mem[16'h04F0] = 8'h00;
mem[16'h04F1] = 8'h08;
mem[16'h04F2] = 8'h18;
mem[16'h04F3] = 8'h3A;
mem[16'h04F4] = 8'h7B;
mem[16'h04F5] = 8'h3E;
mem[16'h04F6] = 8'h1C;
mem[16'h04F7] = 8'h7F;
mem[16'h04F8] = 8'h04;
mem[16'h04F9] = 8'h00;
mem[16'h04FA] = 8'h08;
mem[16'h04FB] = 8'h1C;
mem[16'h04FC] = 8'h1C;
mem[16'h04FD] = 8'h08;
mem[16'h04FE] = 8'h1C;
mem[16'h04FF] = 8'h3E;
mem[16'h0500] = 8'h00;
mem[16'h0501] = 8'h00;
mem[16'h0502] = 8'h00;
mem[16'h0503] = 8'h00;
mem[16'h0504] = 8'h00;
mem[16'h0505] = 8'h00;
mem[16'h0506] = 8'h00;
mem[16'h0507] = 8'h00;
mem[16'h0508] = 8'h10;
mem[16'h0509] = 8'h10;
mem[16'h050A] = 8'h10;
mem[16'h050B] = 8'h10;
mem[16'h050C] = 8'h00;
mem[16'h050D] = 8'h00;
mem[16'h050E] = 8'h10;
mem[16'h050F] = 8'h00;
mem[16'h0510] = 8'h24;
mem[16'h0511] = 8'h24;
mem[16'h0512] = 8'h24;
mem[16'h0513] = 8'h00;
mem[16'h0514] = 8'h00;
mem[16'h0515] = 8'h00;
mem[16'h0516] = 8'h00;
mem[16'h0517] = 8'h00;
mem[16'h0518] = 8'h24;
mem[16'h0519] = 8'h24;
mem[16'h051A] = 8'h7E;
mem[16'h051B] = 8'h24;
mem[16'h051C] = 8'h7E;
mem[16'h051D] = 8'h24;
mem[16'h051E] = 8'h24;
mem[16'h051F] = 8'h00;
mem[16'h0520] = 8'h10;
mem[16'h0521] = 8'h78;
mem[16'h0522] = 8'h14;
mem[16'h0523] = 8'h38;
mem[16'h0524] = 8'h50;
mem[16'h0525] = 8'h3C;
mem[16'h0526] = 8'h10;
mem[16'h0527] = 8'h00;
mem[16'h0528] = 8'h00;
mem[16'h0529] = 8'h46;
mem[16'h052A] = 8'h26;
mem[16'h052B] = 8'h10;
mem[16'h052C] = 8'h08;
mem[16'h052D] = 8'h64;
mem[16'h052E] = 8'h62;
mem[16'h052F] = 8'h00;
mem[16'h0530] = 8'h0C;
mem[16'h0531] = 8'h12;
mem[16'h0532] = 8'h12;
mem[16'h0533] = 8'h0C;
mem[16'h0534] = 8'h52;
mem[16'h0535] = 8'h22;
mem[16'h0536] = 8'h5C;
mem[16'h0537] = 8'h00;
mem[16'h0538] = 8'h20;
mem[16'h0539] = 8'h10;
mem[16'h053A] = 8'h08;
mem[16'h053B] = 8'h00;
mem[16'h053C] = 8'h00;
mem[16'h053D] = 8'h00;
mem[16'h053E] = 8'h00;
mem[16'h053F] = 8'h00;
mem[16'h0540] = 8'h20;
mem[16'h0541] = 8'h10;
mem[16'h0542] = 8'h08;
mem[16'h0543] = 8'h08;
mem[16'h0544] = 8'h08;
mem[16'h0545] = 8'h10;
mem[16'h0546] = 8'h20;
mem[16'h0547] = 8'h00;
mem[16'h0548] = 8'h04;
mem[16'h0549] = 8'h08;
mem[16'h054A] = 8'h10;
mem[16'h054B] = 8'h10;
mem[16'h054C] = 8'h10;
mem[16'h054D] = 8'h08;
mem[16'h054E] = 8'h04;
mem[16'h054F] = 8'h00;
mem[16'h0550] = 8'h10;
mem[16'h0551] = 8'h54;
mem[16'h0552] = 8'h38;
mem[16'h0553] = 8'h7C;
mem[16'h0554] = 8'h38;
mem[16'h0555] = 8'h54;
mem[16'h0556] = 8'h10;
mem[16'h0557] = 8'h00;
mem[16'h0558] = 8'h00;
mem[16'h0559] = 8'h10;
mem[16'h055A] = 8'h10;
mem[16'h055B] = 8'h7C;
mem[16'h055C] = 8'h10;
mem[16'h055D] = 8'h10;
mem[16'h055E] = 8'h00;
mem[16'h055F] = 8'h00;
mem[16'h0560] = 8'h00;
mem[16'h0561] = 8'h00;
mem[16'h0562] = 8'h00;
mem[16'h0563] = 8'h00;
mem[16'h0564] = 8'h00;
mem[16'h0565] = 8'h18;
mem[16'h0566] = 8'h18;
mem[16'h0567] = 8'h0C;
mem[16'h0568] = 8'h00;
mem[16'h0569] = 8'h00;
mem[16'h056A] = 8'h00;
mem[16'h056B] = 8'h7E;
mem[16'h056C] = 8'h00;
mem[16'h056D] = 8'h00;
mem[16'h056E] = 8'h00;
mem[16'h056F] = 8'h00;
mem[16'h0570] = 8'h00;
mem[16'h0571] = 8'h00;
mem[16'h0572] = 8'h00;
mem[16'h0573] = 8'h00;
mem[16'h0574] = 8'h00;
mem[16'h0575] = 8'h18;
mem[16'h0576] = 8'h18;
mem[16'h0577] = 8'h00;
mem[16'h0578] = 8'h28;
mem[16'h0579] = 8'h40;
mem[16'h057A] = 8'h20;
mem[16'h057B] = 8'h10;
mem[16'h057C] = 8'h08;
mem[16'h057D] = 8'h04;
mem[16'h057E] = 8'h02;
mem[16'h057F] = 8'h00;
mem[16'h0580] = 8'h3C;
mem[16'h0581] = 8'h42;
mem[16'h0582] = 8'h42;
mem[16'h0583] = 8'h42;
mem[16'h0584] = 8'h42;
mem[16'h0585] = 8'h42;
mem[16'h0586] = 8'h3C;
mem[16'h0587] = 8'h00;
mem[16'h0588] = 8'h10;
mem[16'h0589] = 8'h18;
mem[16'h058A] = 8'h14;
mem[16'h058B] = 8'h10;
mem[16'h058C] = 8'h10;
mem[16'h058D] = 8'h10;
mem[16'h058E] = 8'h7C;
mem[16'h058F] = 8'h00;
mem[16'h0590] = 8'h3C;
mem[16'h0591] = 8'h42;
mem[16'h0592] = 8'h40;
mem[16'h0593] = 8'h30;
mem[16'h0594] = 8'h0C;
mem[16'h0595] = 8'h02;
mem[16'h0596] = 8'h7E;
mem[16'h0597] = 8'h00;
mem[16'h0598] = 8'h3C;
mem[16'h0599] = 8'h42;
mem[16'h059A] = 8'h40;
mem[16'h059B] = 8'h38;
mem[16'h059C] = 8'h40;
mem[16'h059D] = 8'h42;
mem[16'h059E] = 8'h3C;
mem[16'h059F] = 8'h00;
mem[16'h05A0] = 8'h20;
mem[16'h05A1] = 8'h30;
mem[16'h05A2] = 8'h28;
mem[16'h05A3] = 8'h24;
mem[16'h05A4] = 8'h7E;
mem[16'h05A5] = 8'h20;
mem[16'h05A6] = 8'h20;
mem[16'h05A7] = 8'h00;
mem[16'h05A8] = 8'h7E;
mem[16'h05A9] = 8'h02;
mem[16'h05AA] = 8'h1E;
mem[16'h05AB] = 8'h20;
mem[16'h05AC] = 8'h40;
mem[16'h05AD] = 8'h22;
mem[16'h05AE] = 8'h1C;
mem[16'h05AF] = 8'h00;
mem[16'h05B0] = 8'h38;
mem[16'h05B1] = 8'h04;
mem[16'h05B2] = 8'h02;
mem[16'h05B3] = 8'h3E;
mem[16'h05B4] = 8'h42;
mem[16'h05B5] = 8'h42;
mem[16'h05B6] = 8'h3C;
mem[16'h05B7] = 8'h00;
mem[16'h05B8] = 8'h7E;
mem[16'h05B9] = 8'h42;
mem[16'h05BA] = 8'h20;
mem[16'h05BB] = 8'h10;
mem[16'h05BC] = 8'h08;
mem[16'h05BD] = 8'h08;
mem[16'h05BE] = 8'h08;
mem[16'h05BF] = 8'h00;
mem[16'h05C0] = 8'h3C;
mem[16'h05C1] = 8'h42;
mem[16'h05C2] = 8'h42;
mem[16'h05C3] = 8'h3C;
mem[16'h05C4] = 8'h42;
mem[16'h05C5] = 8'h42;
mem[16'h05C6] = 8'h3C;
mem[16'h05C7] = 8'h00;
mem[16'h05C8] = 8'h3C;
mem[16'h05C9] = 8'h42;
mem[16'h05CA] = 8'h42;
mem[16'h05CB] = 8'h7C;
mem[16'h05CC] = 8'h40;
mem[16'h05CD] = 8'h20;
mem[16'h05CE] = 8'h1C;
mem[16'h05CF] = 8'h00;
mem[16'h05D0] = 8'h00;
mem[16'h05D1] = 8'h00;
mem[16'h05D2] = 8'h18;
mem[16'h05D3] = 8'h18;
mem[16'h05D4] = 8'h00;
mem[16'h05D5] = 8'h18;
mem[16'h05D6] = 8'h18;
mem[16'h05D7] = 8'h00;
mem[16'h05D8] = 8'h00;
mem[16'h05D9] = 8'h00;
mem[16'h05DA] = 8'h18;
mem[16'h05DB] = 8'h18;
mem[16'h05DC] = 8'h00;
mem[16'h05DD] = 8'h18;
mem[16'h05DE] = 8'h18;
mem[16'h05DF] = 8'h0C;
mem[16'h05E0] = 8'h20;
mem[16'h05E1] = 8'h10;
mem[16'h05E2] = 8'h08;
mem[16'h05E3] = 8'h04;
mem[16'h05E4] = 8'h08;
mem[16'h05E5] = 8'h10;
mem[16'h05E6] = 8'h20;
mem[16'h05E7] = 8'h00;
mem[16'h05E8] = 8'h00;
mem[16'h05E9] = 8'h00;
mem[16'h05EA] = 8'h3E;
mem[16'h05EB] = 8'h00;
mem[16'h05EC] = 8'h3E;
mem[16'h05ED] = 8'h00;
mem[16'h05EE] = 8'h00;
mem[16'h05EF] = 8'h00;
mem[16'h05F0] = 8'h04;
mem[16'h05F1] = 8'h08;
mem[16'h05F2] = 8'h10;
mem[16'h05F3] = 8'h20;
mem[16'h05F4] = 8'h10;
mem[16'h05F5] = 8'h08;
mem[16'h05F6] = 8'h04;
mem[16'h05F7] = 8'h00;
mem[16'h05F8] = 8'h60;
mem[16'h05F9] = 8'h42;
mem[16'h05FA] = 8'h40;
mem[16'h05FB] = 8'h30;
mem[16'h05FC] = 8'h08;
mem[16'h05FD] = 8'h00;
mem[16'h05FE] = 8'h08;
mem[16'h05FF] = 8'h00;
mem[16'h0600] = 8'h38;
mem[16'h0601] = 8'h44;
mem[16'h0602] = 8'h52;
mem[16'h0603] = 8'h6A;
mem[16'h0604] = 8'h32;
mem[16'h0605] = 8'h04;
mem[16'h0606] = 8'h78;
mem[16'h0607] = 8'h00;
mem[16'h0608] = 8'h18;
mem[16'h0609] = 8'h24;
mem[16'h060A] = 8'h42;
mem[16'h060B] = 8'h7E;
mem[16'h060C] = 8'h42;
mem[16'h060D] = 8'h42;
mem[16'h060E] = 8'h42;
mem[16'h060F] = 8'h00;
mem[16'h0610] = 8'h3E;
mem[16'h0611] = 8'h44;
mem[16'h0612] = 8'h44;
mem[16'h0613] = 8'h3C;
mem[16'h0614] = 8'h44;
mem[16'h0615] = 8'h44;
mem[16'h0616] = 8'h3E;
mem[16'h0617] = 8'h00;
mem[16'h0618] = 8'h3C;
mem[16'h0619] = 8'h42;
mem[16'h061A] = 8'h02;
mem[16'h061B] = 8'h02;
mem[16'h061C] = 8'h02;
mem[16'h061D] = 8'h42;
mem[16'h061E] = 8'h3C;
mem[16'h061F] = 8'h00;
mem[16'h0620] = 8'h3E;
mem[16'h0621] = 8'h44;
mem[16'h0622] = 8'h44;
mem[16'h0623] = 8'h44;
mem[16'h0624] = 8'h44;
mem[16'h0625] = 8'h44;
mem[16'h0626] = 8'h3E;
mem[16'h0627] = 8'h00;
mem[16'h0628] = 8'h7E;
mem[16'h0629] = 8'h02;
mem[16'h062A] = 8'h02;
mem[16'h062B] = 8'h1E;
mem[16'h062C] = 8'h02;
mem[16'h062D] = 8'h02;
mem[16'h062E] = 8'h7E;
mem[16'h062F] = 8'h00;
mem[16'h0630] = 8'h7E;
mem[16'h0631] = 8'h02;
mem[16'h0632] = 8'h02;
mem[16'h0633] = 8'h1E;
mem[16'h0634] = 8'h02;
mem[16'h0635] = 8'h02;
mem[16'h0636] = 8'h02;
mem[16'h0637] = 8'h00;
mem[16'h0638] = 8'h3C;
mem[16'h0639] = 8'h42;
mem[16'h063A] = 8'h02;
mem[16'h063B] = 8'h72;
mem[16'h063C] = 8'h42;
mem[16'h063D] = 8'h42;
mem[16'h063E] = 8'h3C;
mem[16'h063F] = 8'h00;
mem[16'h0640] = 8'h42;
mem[16'h0641] = 8'h42;
mem[16'h0642] = 8'h42;
mem[16'h0643] = 8'h7E;
mem[16'h0644] = 8'h42;
mem[16'h0645] = 8'h42;
mem[16'h0646] = 8'h42;
mem[16'h0647] = 8'h00;
mem[16'h0648] = 8'h38;
mem[16'h0649] = 8'h10;
mem[16'h064A] = 8'h10;
mem[16'h064B] = 8'h10;
mem[16'h064C] = 8'h10;
mem[16'h064D] = 8'h10;
mem[16'h064E] = 8'h38;
mem[16'h064F] = 8'h00;
mem[16'h0650] = 8'h70;
mem[16'h0651] = 8'h20;
mem[16'h0652] = 8'h20;
mem[16'h0653] = 8'h20;
mem[16'h0654] = 8'h20;
mem[16'h0655] = 8'h22;
mem[16'h0656] = 8'h1C;
mem[16'h0657] = 8'h00;
mem[16'h0658] = 8'h42;
mem[16'h0659] = 8'h22;
mem[16'h065A] = 8'h12;
mem[16'h065B] = 8'h0E;
mem[16'h065C] = 8'h12;
mem[16'h065D] = 8'h22;
mem[16'h065E] = 8'h42;
mem[16'h065F] = 8'h00;
mem[16'h0660] = 8'h02;
mem[16'h0661] = 8'h02;
mem[16'h0662] = 8'h02;
mem[16'h0663] = 8'h02;
mem[16'h0664] = 8'h02;
mem[16'h0665] = 8'h02;
mem[16'h0666] = 8'h7E;
mem[16'h0667] = 8'h00;
mem[16'h0668] = 8'h42;
mem[16'h0669] = 8'h66;
mem[16'h066A] = 8'h5A;
mem[16'h066B] = 8'h5A;
mem[16'h066C] = 8'h42;
mem[16'h066D] = 8'h42;
mem[16'h066E] = 8'h42;
mem[16'h066F] = 8'h00;
mem[16'h0670] = 8'h42;
mem[16'h0671] = 8'h46;
mem[16'h0672] = 8'h4A;
mem[16'h0673] = 8'h52;
mem[16'h0674] = 8'h62;
mem[16'h0675] = 8'h42;
mem[16'h0676] = 8'h42;
mem[16'h0677] = 8'h00;
mem[16'h0678] = 8'h3C;
mem[16'h0679] = 8'h42;
mem[16'h067A] = 8'h42;
mem[16'h067B] = 8'h42;
mem[16'h067C] = 8'h42;
mem[16'h067D] = 8'h42;
mem[16'h067E] = 8'h3C;
mem[16'h067F] = 8'h00;
mem[16'h0680] = 8'h3E;
mem[16'h0681] = 8'h42;
mem[16'h0682] = 8'h42;
mem[16'h0683] = 8'h3E;
mem[16'h0684] = 8'h02;
mem[16'h0685] = 8'h02;
mem[16'h0686] = 8'h02;
mem[16'h0687] = 8'h00;
mem[16'h0688] = 8'h3C;
mem[16'h0689] = 8'h42;
mem[16'h068A] = 8'h42;
mem[16'h068B] = 8'h42;
mem[16'h068C] = 8'h52;
mem[16'h068D] = 8'h22;
mem[16'h068E] = 8'h5C;
mem[16'h068F] = 8'h00;
mem[16'h0690] = 8'h3E;
mem[16'h0691] = 8'h42;
mem[16'h0692] = 8'h42;
mem[16'h0693] = 8'h3E;
mem[16'h0694] = 8'h12;
mem[16'h0695] = 8'h22;
mem[16'h0696] = 8'h42;
mem[16'h0697] = 8'h00;
mem[16'h0698] = 8'h3C;
mem[16'h0699] = 8'h42;
mem[16'h069A] = 8'h02;
mem[16'h069B] = 8'h3C;
mem[16'h069C] = 8'h40;
mem[16'h069D] = 8'h42;
mem[16'h069E] = 8'h3C;
mem[16'h069F] = 8'h00;
mem[16'h06A0] = 8'h7C;
mem[16'h06A1] = 8'h10;
mem[16'h06A2] = 8'h10;
mem[16'h06A3] = 8'h10;
mem[16'h06A4] = 8'h10;
mem[16'h06A5] = 8'h10;
mem[16'h06A6] = 8'h10;
mem[16'h06A7] = 8'h00;
mem[16'h06A8] = 8'h42;
mem[16'h06A9] = 8'h42;
mem[16'h06AA] = 8'h42;
mem[16'h06AB] = 8'h42;
mem[16'h06AC] = 8'h42;
mem[16'h06AD] = 8'h42;
mem[16'h06AE] = 8'h3C;
mem[16'h06AF] = 8'h00;
mem[16'h06B0] = 8'h42;
mem[16'h06B1] = 8'h42;
mem[16'h06B2] = 8'h42;
mem[16'h06B3] = 8'h24;
mem[16'h06B4] = 8'h24;
mem[16'h06B5] = 8'h18;
mem[16'h06B6] = 8'h18;
mem[16'h06B7] = 8'h00;
mem[16'h06B8] = 8'h42;
mem[16'h06B9] = 8'h42;
mem[16'h06BA] = 8'h42;
mem[16'h06BB] = 8'h5A;
mem[16'h06BC] = 8'h5A;
mem[16'h06BD] = 8'h66;
mem[16'h06BE] = 8'h42;
mem[16'h06BF] = 8'h00;
mem[16'h06C0] = 8'h42;
mem[16'h06C1] = 8'h42;
mem[16'h06C2] = 8'h24;
mem[16'h06C3] = 8'h18;
mem[16'h06C4] = 8'h24;
mem[16'h06C5] = 8'h42;
mem[16'h06C6] = 8'h42;
mem[16'h06C7] = 8'h00;
mem[16'h06C8] = 8'h44;
mem[16'h06C9] = 8'h44;
mem[16'h06CA] = 8'h44;
mem[16'h06CB] = 8'h38;
mem[16'h06CC] = 8'h10;
mem[16'h06CD] = 8'h10;
mem[16'h06CE] = 8'h10;
mem[16'h06CF] = 8'h00;
mem[16'h06D0] = 8'h7E;
mem[16'h06D1] = 8'h40;
mem[16'h06D2] = 8'h20;
mem[16'h06D3] = 8'h18;
mem[16'h06D4] = 8'h04;
mem[16'h06D5] = 8'h02;
mem[16'h06D6] = 8'h7E;
mem[16'h06D7] = 8'h00;
mem[16'h06D8] = 8'h3C;
mem[16'h06D9] = 8'h04;
mem[16'h06DA] = 8'h04;
mem[16'h06DB] = 8'h04;
mem[16'h06DC] = 8'h04;
mem[16'h06DD] = 8'h04;
mem[16'h06DE] = 8'h3C;
mem[16'h06DF] = 8'h00;
mem[16'h06E0] = 8'h00;
mem[16'h06E1] = 8'h02;
mem[16'h06E2] = 8'h04;
mem[16'h06E3] = 8'h08;
mem[16'h06E4] = 8'h10;
mem[16'h06E5] = 8'h20;
mem[16'h06E6] = 8'h40;
mem[16'h06E7] = 8'h00;
mem[16'h06E8] = 8'h3C;
mem[16'h06E9] = 8'h20;
mem[16'h06EA] = 8'h20;
mem[16'h06EB] = 8'h20;
mem[16'h06EC] = 8'h20;
mem[16'h06ED] = 8'h20;
mem[16'h06EE] = 8'h3C;
mem[16'h06EF] = 8'h00;
mem[16'h06F0] = 8'h10;
mem[16'h06F1] = 8'h28;
mem[16'h06F2] = 8'h44;
mem[16'h06F3] = 8'h00;
mem[16'h06F4] = 8'h00;
mem[16'h06F5] = 8'h00;
mem[16'h06F6] = 8'h00;
mem[16'h06F7] = 8'h00;
mem[16'h06F8] = 8'h02;
mem[16'h06F9] = 8'h00;
mem[16'h06FA] = 8'h00;
mem[16'h06FB] = 8'h00;
mem[16'h06FC] = 8'h00;
mem[16'h06FD] = 8'h00;
mem[16'h06FE] = 8'h00;
mem[16'h06FF] = 8'hFF;
mem[16'h0700] = 8'h08;
mem[16'h0701] = 8'h10;
mem[16'h0702] = 8'h20;
mem[16'h0703] = 8'h00;
mem[16'h0704] = 8'h00;
mem[16'h0705] = 8'h00;
mem[16'h0706] = 8'h00;
mem[16'h0707] = 8'h00;
mem[16'h0708] = 8'h00;
mem[16'h0709] = 8'h00;
mem[16'h070A] = 8'h1C;
mem[16'h070B] = 8'h20;
mem[16'h070C] = 8'h3C;
mem[16'h070D] = 8'h22;
mem[16'h070E] = 8'h5C;
mem[16'h070F] = 8'h00;
mem[16'h0710] = 8'h02;
mem[16'h0711] = 8'h02;
mem[16'h0712] = 8'h3A;
mem[16'h0713] = 8'h46;
mem[16'h0714] = 8'h42;
mem[16'h0715] = 8'h46;
mem[16'h0716] = 8'h3A;
mem[16'h0717] = 8'h00;
mem[16'h0718] = 8'h00;
mem[16'h0719] = 8'h00;
mem[16'h071A] = 8'h3C;
mem[16'h071B] = 8'h02;
mem[16'h071C] = 8'h02;
mem[16'h071D] = 8'h02;
mem[16'h071E] = 8'h3C;
mem[16'h071F] = 8'h00;
mem[16'h0720] = 8'h40;
mem[16'h0721] = 8'h40;
mem[16'h0722] = 8'h5C;
mem[16'h0723] = 8'h62;
mem[16'h0724] = 8'h42;
mem[16'h0725] = 8'h62;
mem[16'h0726] = 8'h5C;
mem[16'h0727] = 8'h00;
mem[16'h0728] = 8'h00;
mem[16'h0729] = 8'h00;
mem[16'h072A] = 8'h3C;
mem[16'h072B] = 8'h42;
mem[16'h072C] = 8'h7E;
mem[16'h072D] = 8'h02;
mem[16'h072E] = 8'h3C;
mem[16'h072F] = 8'h00;
mem[16'h0730] = 8'h30;
mem[16'h0731] = 8'h48;
mem[16'h0732] = 8'h08;
mem[16'h0733] = 8'h3E;
mem[16'h0734] = 8'h08;
mem[16'h0735] = 8'h08;
mem[16'h0736] = 8'h08;
mem[16'h0737] = 8'h00;
mem[16'h0738] = 8'h00;
mem[16'h0739] = 8'h00;
mem[16'h073A] = 8'h5C;
mem[16'h073B] = 8'h62;
mem[16'h073C] = 8'h62;
mem[16'h073D] = 8'h5C;
mem[16'h073E] = 8'h40;
mem[16'h073F] = 8'h3C;
mem[16'h0740] = 8'h02;
mem[16'h0741] = 8'h02;
mem[16'h0742] = 8'h3A;
mem[16'h0743] = 8'h46;
mem[16'h0744] = 8'h42;
mem[16'h0745] = 8'h42;
mem[16'h0746] = 8'h42;
mem[16'h0747] = 8'h00;
mem[16'h0748] = 8'h10;
mem[16'h0749] = 8'h00;
mem[16'h074A] = 8'h18;
mem[16'h074B] = 8'h10;
mem[16'h074C] = 8'h10;
mem[16'h074D] = 8'h10;
mem[16'h074E] = 8'h38;
mem[16'h074F] = 8'h00;
mem[16'h0750] = 8'h20;
mem[16'h0751] = 8'h00;
mem[16'h0752] = 8'h30;
mem[16'h0753] = 8'h20;
mem[16'h0754] = 8'h20;
mem[16'h0755] = 8'h20;
mem[16'h0756] = 8'h22;
mem[16'h0757] = 8'h1C;
mem[16'h0758] = 8'h02;
mem[16'h0759] = 8'h02;
mem[16'h075A] = 8'h22;
mem[16'h075B] = 8'h12;
mem[16'h075C] = 8'h0A;
mem[16'h075D] = 8'h16;
mem[16'h075E] = 8'h22;
mem[16'h075F] = 8'h00;
mem[16'h0760] = 8'h18;
mem[16'h0761] = 8'h10;
mem[16'h0762] = 8'h10;
mem[16'h0763] = 8'h10;
mem[16'h0764] = 8'h10;
mem[16'h0765] = 8'h10;
mem[16'h0766] = 8'h38;
mem[16'h0767] = 8'h00;
mem[16'h0768] = 8'h00;
mem[16'h0769] = 8'h00;
mem[16'h076A] = 8'h2E;
mem[16'h076B] = 8'h54;
mem[16'h076C] = 8'h54;
mem[16'h076D] = 8'h54;
mem[16'h076E] = 8'h54;
mem[16'h076F] = 8'h00;
mem[16'h0770] = 8'h00;
mem[16'h0771] = 8'h00;
mem[16'h0772] = 8'h3E;
mem[16'h0773] = 8'h44;
mem[16'h0774] = 8'h44;
mem[16'h0775] = 8'h44;
mem[16'h0776] = 8'h44;
mem[16'h0777] = 8'h00;
mem[16'h0778] = 8'h00;
mem[16'h0779] = 8'h00;
mem[16'h077A] = 8'h38;
mem[16'h077B] = 8'h44;
mem[16'h077C] = 8'h44;
mem[16'h077D] = 8'h44;
mem[16'h077E] = 8'h38;
mem[16'h077F] = 8'h00;
mem[16'h0780] = 8'h00;
mem[16'h0781] = 8'h00;
mem[16'h0782] = 8'h3A;
mem[16'h0783] = 8'h46;
mem[16'h0784] = 8'h46;
mem[16'h0785] = 8'h3A;
mem[16'h0786] = 8'h02;
mem[16'h0787] = 8'h02;
mem[16'h0788] = 8'h00;
mem[16'h0789] = 8'h00;
mem[16'h078A] = 8'h5C;
mem[16'h078B] = 8'h62;
mem[16'h078C] = 8'h62;
mem[16'h078D] = 8'h5C;
mem[16'h078E] = 8'h40;
mem[16'h078F] = 8'h40;
mem[16'h0790] = 8'h00;
mem[16'h0791] = 8'h00;
mem[16'h0792] = 8'h3A;
mem[16'h0793] = 8'h46;
mem[16'h0794] = 8'h02;
mem[16'h0795] = 8'h02;
mem[16'h0796] = 8'h02;
mem[16'h0797] = 8'h00;
mem[16'h0798] = 8'h00;
mem[16'h0799] = 8'h00;
mem[16'h079A] = 8'h7C;
mem[16'h079B] = 8'h02;
mem[16'h079C] = 8'h3C;
mem[16'h079D] = 8'h40;
mem[16'h079E] = 8'h3E;
mem[16'h079F] = 8'h00;
mem[16'h07A0] = 8'h08;
mem[16'h07A1] = 8'h08;
mem[16'h07A2] = 8'h3E;
mem[16'h07A3] = 8'h08;
mem[16'h07A4] = 8'h08;
mem[16'h07A5] = 8'h48;
mem[16'h07A6] = 8'h30;
mem[16'h07A7] = 8'h00;
mem[16'h07A8] = 8'h00;
mem[16'h07A9] = 8'h00;
mem[16'h07AA] = 8'h42;
mem[16'h07AB] = 8'h42;
mem[16'h07AC] = 8'h42;
mem[16'h07AD] = 8'h62;
mem[16'h07AE] = 8'h5C;
mem[16'h07AF] = 8'h00;
mem[16'h07B0] = 8'h00;
mem[16'h07B1] = 8'h00;
mem[16'h07B2] = 8'h42;
mem[16'h07B3] = 8'h42;
mem[16'h07B4] = 8'h42;
mem[16'h07B5] = 8'h24;
mem[16'h07B6] = 8'h18;
mem[16'h07B7] = 8'h00;
mem[16'h07B8] = 8'h00;
mem[16'h07B9] = 8'h00;
mem[16'h07BA] = 8'h44;
mem[16'h07BB] = 8'h44;
mem[16'h07BC] = 8'h54;
mem[16'h07BD] = 8'h54;
mem[16'h07BE] = 8'h6C;
mem[16'h07BF] = 8'h00;
mem[16'h07C0] = 8'h00;
mem[16'h07C1] = 8'h00;
mem[16'h07C2] = 8'h42;
mem[16'h07C3] = 8'h24;
mem[16'h07C4] = 8'h18;
mem[16'h07C5] = 8'h24;
mem[16'h07C6] = 8'h42;
mem[16'h07C7] = 8'h00;
mem[16'h07C8] = 8'h00;
mem[16'h07C9] = 8'h00;
mem[16'h07CA] = 8'h42;
mem[16'h07CB] = 8'h42;
mem[16'h07CC] = 8'h62;
mem[16'h07CD] = 8'h5C;
mem[16'h07CE] = 8'h40;
mem[16'h07CF] = 8'h3C;
mem[16'h07D0] = 8'h00;
mem[16'h07D1] = 8'h00;
mem[16'h07D2] = 8'h7E;
mem[16'h07D3] = 8'h20;
mem[16'h07D4] = 8'h18;
mem[16'h07D5] = 8'h04;
mem[16'h07D6] = 8'h7E;
mem[16'h07D7] = 8'h00;
mem[16'h07D8] = 8'h38;
mem[16'h07D9] = 8'h04;
mem[16'h07DA] = 8'h04;
mem[16'h07DB] = 8'h06;
mem[16'h07DC] = 8'h04;
mem[16'h07DD] = 8'h04;
mem[16'h07DE] = 8'h38;
mem[16'h07DF] = 8'h00;
mem[16'h07E0] = 8'h08;
mem[16'h07E1] = 8'h08;
mem[16'h07E2] = 8'h08;
mem[16'h07E3] = 8'h08;
mem[16'h07E4] = 8'h08;
mem[16'h07E5] = 8'h08;
mem[16'h07E6] = 8'h08;
mem[16'h07E7] = 8'h08;
mem[16'h07E8] = 8'h0E;
mem[16'h07E9] = 8'h10;
mem[16'h07EA] = 8'h10;
mem[16'h07EB] = 8'h30;
mem[16'h07EC] = 8'h10;
mem[16'h07ED] = 8'h10;
mem[16'h07EE] = 8'h0E;
mem[16'h07EF] = 8'h00;
mem[16'h07F0] = 8'h28;
mem[16'h07F1] = 8'h14;
mem[16'h07F2] = 8'h00;
mem[16'h07F3] = 8'h00;
mem[16'h07F4] = 8'h00;
mem[16'h07F5] = 8'h00;
mem[16'h07F6] = 8'h00;
mem[16'h07F7] = 8'h00;
mem[16'h07F8] = 8'hFF;
mem[16'h07F9] = 8'hFF;
mem[16'h07FA] = 8'hFF;
mem[16'h07FB] = 8'hFF;
mem[16'h07FC] = 8'hFF;
mem[16'h07FD] = 8'h0F;
mem[16'h07FE] = 8'hAB;
mem[16'h07FF] = 8'h81;
mem[16'h0800] = 8'h4C;
mem[16'h0801] = 8'h00;
mem[16'h0802] = 8'h0C;
mem[16'h0803] = 8'hAA;
mem[16'h0804] = 8'hAA;
mem[16'h0805] = 8'hAA;
mem[16'h0806] = 8'hAA;
mem[16'h0807] = 8'hAA;
mem[16'h0808] = 8'hAA;
mem[16'h0809] = 8'hAA;
mem[16'h080A] = 8'hAA;
mem[16'h080B] = 8'hAA;
mem[16'h080C] = 8'hAA;
mem[16'h080D] = 8'hAA;
mem[16'h080E] = 8'hAA;
mem[16'h080F] = 8'hAA;
mem[16'h0810] = 8'hAA;
mem[16'h0811] = 8'hAA;
mem[16'h0812] = 8'hAA;
mem[16'h0813] = 8'hAA;
mem[16'h0814] = 8'hAA;
mem[16'h0815] = 8'hAA;
mem[16'h0816] = 8'hAA;
mem[16'h0817] = 8'hAA;
mem[16'h0818] = 8'hAA;
mem[16'h0819] = 8'hAA;
mem[16'h081A] = 8'hAA;
mem[16'h081B] = 8'hAA;
mem[16'h081C] = 8'hAA;
mem[16'h081D] = 8'hAA;
mem[16'h081E] = 8'hAA;
mem[16'h081F] = 8'hAA;
mem[16'h0820] = 8'hAA;
mem[16'h0821] = 8'hAA;
mem[16'h0822] = 8'hAA;
mem[16'h0823] = 8'hAA;
mem[16'h0824] = 8'hAA;
mem[16'h0825] = 8'hAA;
mem[16'h0826] = 8'hAA;
mem[16'h0827] = 8'hA0;
mem[16'h0828] = 8'hAA;
mem[16'h0829] = 8'hAA;
mem[16'h082A] = 8'hA0;
mem[16'h082B] = 8'hA0;
mem[16'h082C] = 8'hA0;
mem[16'h082D] = 8'hA0;
mem[16'h082E] = 8'hA0;
mem[16'h082F] = 8'hA0;
mem[16'h0830] = 8'hA0;
mem[16'h0831] = 8'hA0;
mem[16'h0832] = 8'hA0;
mem[16'h0833] = 8'hA0;
mem[16'h0834] = 8'hA0;
mem[16'h0835] = 8'hA0;
mem[16'h0836] = 8'hA0;
mem[16'h0837] = 8'hA0;
mem[16'h0838] = 8'hA0;
mem[16'h0839] = 8'hA0;
mem[16'h083A] = 8'hA0;
mem[16'h083B] = 8'hA0;
mem[16'h083C] = 8'hA0;
mem[16'h083D] = 8'hA0;
mem[16'h083E] = 8'hA0;
mem[16'h083F] = 8'hA0;
mem[16'h0840] = 8'hA0;
mem[16'h0841] = 8'hA0;
mem[16'h0842] = 8'hA0;
mem[16'h0843] = 8'hA0;
mem[16'h0844] = 8'hA0;
mem[16'h0845] = 8'hA0;
mem[16'h0846] = 8'hA0;
mem[16'h0847] = 8'hA0;
mem[16'h0848] = 8'hA0;
mem[16'h0849] = 8'hA0;
mem[16'h084A] = 8'hA0;
mem[16'h084B] = 8'hA0;
mem[16'h084C] = 8'hA0;
mem[16'h084D] = 8'hAA;
mem[16'h084E] = 8'hAA;
mem[16'h084F] = 8'hA0;
mem[16'h0850] = 8'hAA;
mem[16'h0851] = 8'hAA;
mem[16'h0852] = 8'hA0;
mem[16'h0853] = 8'hA0;
mem[16'h0854] = 8'hA0;
mem[16'h0855] = 8'hA0;
mem[16'h0856] = 8'hA0;
mem[16'h0857] = 8'hA0;
mem[16'h0858] = 8'hA0;
mem[16'h0859] = 8'hA0;
mem[16'h085A] = 8'hA0;
mem[16'h085B] = 8'hA0;
mem[16'h085C] = 8'hA0;
mem[16'h085D] = 8'hA0;
mem[16'h085E] = 8'hA0;
mem[16'h085F] = 8'hA0;
mem[16'h0860] = 8'hA0;
mem[16'h0861] = 8'hA0;
mem[16'h0862] = 8'hA0;
mem[16'h0863] = 8'hA0;
mem[16'h0864] = 8'hA0;
mem[16'h0865] = 8'hA0;
mem[16'h0866] = 8'hA0;
mem[16'h0867] = 8'hA0;
mem[16'h0868] = 8'hA0;
mem[16'h0869] = 8'hA0;
mem[16'h086A] = 8'hA0;
mem[16'h086B] = 8'hA0;
mem[16'h086C] = 8'hA0;
mem[16'h086D] = 8'hA0;
mem[16'h086E] = 8'hA0;
mem[16'h086F] = 8'hA0;
mem[16'h0870] = 8'hA0;
mem[16'h0871] = 8'hA0;
mem[16'h0872] = 8'hA0;
mem[16'h0873] = 8'hA0;
mem[16'h0874] = 8'hA0;
mem[16'h0875] = 8'hAA;
mem[16'h0876] = 8'hAA;
mem[16'h0877] = 8'hA0;
mem[16'h0878] = 8'h1D;
mem[16'h0879] = 8'h00;
mem[16'h087A] = 8'h00;
mem[16'h087B] = 8'h7C;
mem[16'h087C] = 8'h2A;
mem[16'h087D] = 8'h28;
mem[16'h087E] = 8'h3A;
mem[16'h087F] = 8'h00;
mem[16'h0880] = 8'hAA;
mem[16'h0881] = 8'hAA;
mem[16'h0882] = 8'hAA;
mem[16'h0883] = 8'hA0;
mem[16'h0884] = 8'hA0;
mem[16'h0885] = 8'hA0;
mem[16'h0886] = 8'hA0;
mem[16'h0887] = 8'hA0;
mem[16'h0888] = 8'hA0;
mem[16'h0889] = 8'hA0;
mem[16'h088A] = 8'hA0;
mem[16'h088B] = 8'hA0;
mem[16'h088C] = 8'hA0;
mem[16'h088D] = 8'hA0;
mem[16'h088E] = 8'hA0;
mem[16'h088F] = 8'hA0;
mem[16'h0890] = 8'hA0;
mem[16'h0891] = 8'hA0;
mem[16'h0892] = 8'hA0;
mem[16'h0893] = 8'hA0;
mem[16'h0894] = 8'hA0;
mem[16'h0895] = 8'hA0;
mem[16'h0896] = 8'hA0;
mem[16'h0897] = 8'hA0;
mem[16'h0898] = 8'hA0;
mem[16'h0899] = 8'hA0;
mem[16'h089A] = 8'hA0;
mem[16'h089B] = 8'hA0;
mem[16'h089C] = 8'hA0;
mem[16'h089D] = 8'hA0;
mem[16'h089E] = 8'hA0;
mem[16'h089F] = 8'hA0;
mem[16'h08A0] = 8'hA0;
mem[16'h08A1] = 8'hA0;
mem[16'h08A2] = 8'hA0;
mem[16'h08A3] = 8'hA0;
mem[16'h08A4] = 8'hAA;
mem[16'h08A5] = 8'hAA;
mem[16'h08A6] = 8'hAA;
mem[16'h08A7] = 8'hA0;
mem[16'h08A8] = 8'hAA;
mem[16'h08A9] = 8'hAA;
mem[16'h08AA] = 8'hA0;
mem[16'h08AB] = 8'hA0;
mem[16'h08AC] = 8'hA0;
mem[16'h08AD] = 8'hA0;
mem[16'h08AE] = 8'hA0;
mem[16'h08AF] = 8'hA0;
mem[16'h08B0] = 8'hA0;
mem[16'h08B1] = 8'hA0;
mem[16'h08B2] = 8'hA0;
mem[16'h08B3] = 8'hA0;
mem[16'h08B4] = 8'hA0;
mem[16'h08B5] = 8'hA0;
mem[16'h08B6] = 8'hA0;
mem[16'h08B7] = 8'hA0;
mem[16'h08B8] = 8'hA0;
mem[16'h08B9] = 8'hA0;
mem[16'h08BA] = 8'hC1;
mem[16'h08BB] = 8'hA0;
mem[16'h08BC] = 8'hA0;
mem[16'h08BD] = 8'hA0;
mem[16'h08BE] = 8'hA0;
mem[16'h08BF] = 8'hA0;
mem[16'h08C0] = 8'hA0;
mem[16'h08C1] = 8'hA0;
mem[16'h08C2] = 8'hA0;
mem[16'h08C3] = 8'hA0;
mem[16'h08C4] = 8'hA0;
mem[16'h08C5] = 8'hA0;
mem[16'h08C6] = 8'hA0;
mem[16'h08C7] = 8'hA0;
mem[16'h08C8] = 8'hA0;
mem[16'h08C9] = 8'hA0;
mem[16'h08CA] = 8'hA0;
mem[16'h08CB] = 8'hA0;
mem[16'h08CC] = 8'hA0;
mem[16'h08CD] = 8'hAA;
mem[16'h08CE] = 8'hAA;
mem[16'h08CF] = 8'hA0;
mem[16'h08D0] = 8'hAA;
mem[16'h08D1] = 8'hAA;
mem[16'h08D2] = 8'hA0;
mem[16'h08D3] = 8'hA0;
mem[16'h08D4] = 8'h0A;
mem[16'h08D5] = 8'hA0;
mem[16'h08D6] = 8'hD4;
mem[16'h08D7] = 8'hCF;
mem[16'h08D8] = 8'hA0;
mem[16'h08D9] = 8'hC6;
mem[16'h08DA] = 8'hD2;
mem[16'h08DB] = 8'hCF;
mem[16'h08DC] = 8'hC7;
mem[16'h08DD] = 8'hA0;
mem[16'h08DE] = 8'hD7;
mem[16'h08DF] = 8'hC9;
mem[16'h08E0] = 8'hD4;
mem[16'h08E1] = 8'hC8;
mem[16'h08E2] = 8'hA0;
mem[16'h08E3] = 8'hD9;
mem[16'h08E4] = 8'hCF;
mem[16'h08E5] = 8'hD5;
mem[16'h08E6] = 8'hD2;
mem[16'h08E7] = 8'hA0;
mem[16'h08E8] = 8'hCA;
mem[16'h08E9] = 8'hCF;
mem[16'h08EA] = 8'hD9;
mem[16'h08EB] = 8'hD3;
mem[16'h08EC] = 8'hD4;
mem[16'h08ED] = 8'hC9;
mem[16'h08EE] = 8'hC3;
mem[16'h08EF] = 8'hCB;
mem[16'h08F0] = 8'hA0;
mem[16'h08F1] = 8'hA0;
mem[16'h08F2] = 8'hA0;
mem[16'h08F3] = 8'hA0;
mem[16'h08F4] = 8'hA0;
mem[16'h08F5] = 8'hAA;
mem[16'h08F6] = 8'hAA;
mem[16'h08F7] = 8'hA0;
mem[16'h08F8] = 8'h04;
mem[16'h08F9] = 8'h00;
mem[16'h08FA] = 8'h08;
mem[16'h08FB] = 8'h1C;
mem[16'h08FC] = 8'h1C;
mem[16'h08FD] = 8'h08;
mem[16'h08FE] = 8'h00;
mem[16'h08FF] = 8'h3E;
mem[16'h0900] = 8'hAA;
mem[16'h0901] = 8'hAA;
mem[16'h0902] = 8'hA0;
mem[16'h0903] = 8'hA0;
mem[16'h0904] = 8'hA0;
mem[16'h0905] = 8'hA0;
mem[16'h0906] = 8'hA0;
mem[16'h0907] = 8'hA0;
mem[16'h0908] = 8'hA0;
mem[16'h0909] = 8'hA0;
mem[16'h090A] = 8'hA0;
mem[16'h090B] = 8'hA0;
mem[16'h090C] = 8'hA0;
mem[16'h090D] = 8'hA0;
mem[16'h090E] = 8'hA0;
mem[16'h090F] = 8'hC6;
mem[16'h0910] = 8'hD2;
mem[16'h0911] = 8'hCF;
mem[16'h0912] = 8'hC7;
mem[16'h0913] = 8'hC7;
mem[16'h0914] = 8'hC5;
mem[16'h0915] = 8'hD2;
mem[16'h0916] = 8'hA0;
mem[16'h0917] = 8'hA0;
mem[16'h0918] = 8'hA0;
mem[16'h0919] = 8'hA0;
mem[16'h091A] = 8'hA0;
mem[16'h091B] = 8'hA0;
mem[16'h091C] = 8'hA0;
mem[16'h091D] = 8'hA0;
mem[16'h091E] = 8'hA0;
mem[16'h091F] = 8'hA0;
mem[16'h0920] = 8'hA0;
mem[16'h0921] = 8'hA0;
mem[16'h0922] = 8'hA0;
mem[16'h0923] = 8'hA0;
mem[16'h0924] = 8'hA0;
mem[16'h0925] = 8'hAA;
mem[16'h0926] = 8'hAA;
mem[16'h0927] = 8'hA0;
mem[16'h0928] = 8'hAA;
mem[16'h0929] = 8'hAA;
mem[16'h092A] = 8'hA0;
mem[16'h092B] = 8'hA0;
mem[16'h092C] = 8'hA0;
mem[16'h092D] = 8'hA0;
mem[16'h092E] = 8'hA0;
mem[16'h092F] = 8'hA0;
mem[16'h0930] = 8'hA0;
mem[16'h0931] = 8'hA0;
mem[16'h0932] = 8'hA0;
mem[16'h0933] = 8'hA0;
mem[16'h0934] = 8'hA0;
mem[16'h0935] = 8'hA0;
mem[16'h0936] = 8'hA0;
mem[16'h0937] = 8'hA0;
mem[16'h0938] = 8'hBC;
mem[16'h0939] = 8'hAD;
mem[16'h093A] = 8'hA0;
mem[16'h093B] = 8'hAD;
mem[16'h093C] = 8'hBE;
mem[16'h093D] = 8'hA0;
mem[16'h093E] = 8'hA0;
mem[16'h093F] = 8'hA0;
mem[16'h0940] = 8'hA0;
mem[16'h0941] = 8'hA0;
mem[16'h0942] = 8'hA0;
mem[16'h0943] = 8'hA0;
mem[16'h0944] = 8'hA0;
mem[16'h0945] = 8'hA0;
mem[16'h0946] = 8'hA0;
mem[16'h0947] = 8'hA0;
mem[16'h0948] = 8'hA0;
mem[16'h0949] = 8'hA0;
mem[16'h094A] = 8'hA0;
mem[16'h094B] = 8'hA0;
mem[16'h094C] = 8'hA0;
mem[16'h094D] = 8'hAA;
mem[16'h094E] = 8'hAA;
mem[16'h094F] = 8'hA0;
mem[16'h0950] = 8'hAA;
mem[16'h0951] = 8'hAA;
mem[16'h0952] = 8'hA0;
mem[16'h0953] = 8'hA0;
mem[16'h0954] = 8'hA0;
mem[16'h0955] = 8'hA0;
mem[16'h0956] = 8'hA0;
mem[16'h0957] = 8'hA0;
mem[16'h0958] = 8'hA0;
mem[16'h0959] = 8'hA0;
mem[16'h095A] = 8'hA0;
mem[16'h095B] = 8'hA0;
mem[16'h095C] = 8'hA0;
mem[16'h095D] = 8'hA0;
mem[16'h095E] = 8'hA0;
mem[16'h095F] = 8'hA0;
mem[16'h0960] = 8'hA0;
mem[16'h0961] = 8'hA0;
mem[16'h0962] = 8'hA0;
mem[16'h0963] = 8'hA0;
mem[16'h0964] = 8'hA0;
mem[16'h0965] = 8'hA0;
mem[16'h0966] = 8'hA0;
mem[16'h0967] = 8'hA0;
mem[16'h0968] = 8'hA0;
mem[16'h0969] = 8'hA0;
mem[16'h096A] = 8'hA0;
mem[16'h096B] = 8'hA0;
mem[16'h096C] = 8'hA0;
mem[16'h096D] = 8'hA0;
mem[16'h096E] = 8'hA0;
mem[16'h096F] = 8'hA0;
mem[16'h0970] = 8'hA0;
mem[16'h0971] = 8'hA0;
mem[16'h0972] = 8'hA0;
mem[16'h0973] = 8'hA0;
mem[16'h0974] = 8'hA0;
mem[16'h0975] = 8'hAA;
mem[16'h0976] = 8'hAA;
mem[16'h0977] = 8'hA0;
mem[16'h0978] = 8'h30;
mem[16'h0979] = 8'h40;
mem[16'h097A] = 8'h20;
mem[16'h097B] = 8'h10;
mem[16'h097C] = 8'h08;
mem[16'h097D] = 8'h04;
mem[16'h097E] = 8'h02;
mem[16'h097F] = 8'h00;
mem[16'h0980] = 8'hAA;
mem[16'h0981] = 8'hAA;
mem[16'h0982] = 8'hA0;
mem[16'h0983] = 8'hA0;
mem[16'h0984] = 8'hA0;
mem[16'h0985] = 8'hA0;
mem[16'h0986] = 8'hA0;
mem[16'h0987] = 8'hA0;
mem[16'h0988] = 8'hA0;
mem[16'h0989] = 8'hC6;
mem[16'h098A] = 8'hD2;
mem[16'h098B] = 8'hCF;
mem[16'h098C] = 8'hCD;
mem[16'h098D] = 8'hA0;
mem[16'h098E] = 8'hD3;
mem[16'h098F] = 8'hC9;
mem[16'h0990] = 8'hC5;
mem[16'h0991] = 8'hD2;
mem[16'h0992] = 8'hD2;
mem[16'h0993] = 8'hC1;
mem[16'h0994] = 8'hA0;
mem[16'h0995] = 8'hCF;
mem[16'h0996] = 8'hCE;
mem[16'h0997] = 8'hAD;
mem[16'h0998] = 8'hCC;
mem[16'h0999] = 8'hC9;
mem[16'h099A] = 8'hCE;
mem[16'h099B] = 8'hC5;
mem[16'h099C] = 8'hA0;
mem[16'h099D] = 8'hA0;
mem[16'h099E] = 8'hA0;
mem[16'h099F] = 8'hA0;
mem[16'h09A0] = 8'hA0;
mem[16'h09A1] = 8'hA0;
mem[16'h09A2] = 8'hA0;
mem[16'h09A3] = 8'hA0;
mem[16'h09A4] = 8'hA0;
mem[16'h09A5] = 8'hAA;
mem[16'h09A6] = 8'hAA;
mem[16'h09A7] = 8'hA0;
mem[16'h09A8] = 8'hAA;
mem[16'h09A9] = 8'hAA;
mem[16'h09AA] = 8'hA0;
mem[16'h09AB] = 8'hA0;
mem[16'h09AC] = 8'hA0;
mem[16'h09AD] = 8'hA0;
mem[16'h09AE] = 8'hA0;
mem[16'h09AF] = 8'hA0;
mem[16'h09B0] = 8'hA0;
mem[16'h09B1] = 8'hA0;
mem[16'h09B2] = 8'hA0;
mem[16'h09B3] = 8'hA0;
mem[16'h09B4] = 8'hA0;
mem[16'h09B5] = 8'hA0;
mem[16'h09B6] = 8'hA0;
mem[16'h09B7] = 8'hA0;
mem[16'h09B8] = 8'hA0;
mem[16'h09B9] = 8'hA0;
mem[16'h09BA] = 8'hDA;
mem[16'h09BB] = 8'hA0;
mem[16'h09BC] = 8'hA0;
mem[16'h09BD] = 8'hA0;
mem[16'h09BE] = 8'hA0;
mem[16'h09BF] = 8'hA0;
mem[16'h09C0] = 8'hA0;
mem[16'h09C1] = 8'hA0;
mem[16'h09C2] = 8'hA0;
mem[16'h09C3] = 8'hA0;
mem[16'h09C4] = 8'hA0;
mem[16'h09C5] = 8'hA0;
mem[16'h09C6] = 8'hA0;
mem[16'h09C7] = 8'hA0;
mem[16'h09C8] = 8'hA0;
mem[16'h09C9] = 8'hA0;
mem[16'h09CA] = 8'hA0;
mem[16'h09CB] = 8'hA0;
mem[16'h09CC] = 8'hA0;
mem[16'h09CD] = 8'hAA;
mem[16'h09CE] = 8'hAA;
mem[16'h09CF] = 8'hA0;
mem[16'h09D0] = 8'hAA;
mem[16'h09D1] = 8'hAA;
mem[16'h09D2] = 8'hA0;
mem[16'h09D3] = 8'hA0;
mem[16'h09D4] = 8'h05;
mem[16'h09D5] = 8'h13;
mem[16'h09D6] = 8'h03;
mem[16'h09D7] = 8'hA0;
mem[16'h09D8] = 8'hD4;
mem[16'h09D9] = 8'hCF;
mem[16'h09DA] = 8'hA0;
mem[16'h09DB] = 8'hD3;
mem[16'h09DC] = 8'hD4;
mem[16'h09DD] = 8'hCF;
mem[16'h09DE] = 8'hD0;
mem[16'h09DF] = 8'hA0;
mem[16'h09E0] = 8'hA0;
mem[16'h09E1] = 8'h21;
mem[16'h09E2] = 8'hA0;
mem[16'h09E3] = 8'hD4;
mem[16'h09E4] = 8'hCF;
mem[16'h09E5] = 8'hA0;
mem[16'h09E6] = 8'hD3;
mem[16'h09E7] = 8'hCC;
mem[16'h09E8] = 8'hCF;
mem[16'h09E9] = 8'hD7;
mem[16'h09EA] = 8'hA0;
mem[16'h09EB] = 8'hC7;
mem[16'h09EC] = 8'hC1;
mem[16'h09ED] = 8'hCD;
mem[16'h09EE] = 8'hC5;
mem[16'h09EF] = 8'hA0;
mem[16'h09F0] = 8'hA0;
mem[16'h09F1] = 8'hA0;
mem[16'h09F2] = 8'hA0;
mem[16'h09F3] = 8'hA0;
mem[16'h09F4] = 8'hA0;
mem[16'h09F5] = 8'hAA;
mem[16'h09F6] = 8'hAA;
mem[16'h09F7] = 8'hA0;
mem[16'h09F8] = 8'h60;
mem[16'h09F9] = 8'h42;
mem[16'h09FA] = 8'h40;
mem[16'h09FB] = 8'h30;
mem[16'h09FC] = 8'h08;
mem[16'h09FD] = 8'h00;
mem[16'h09FE] = 8'h08;
mem[16'h09FF] = 8'h00;
mem[16'h0A00] = 8'hAA;
mem[16'h0A01] = 8'hAA;
mem[16'h0A02] = 8'hA0;
mem[16'h0A03] = 8'hA0;
mem[16'h0A04] = 8'hA0;
mem[16'h0A05] = 8'hA0;
mem[16'h0A06] = 8'hA0;
mem[16'h0A07] = 8'hA0;
mem[16'h0A08] = 8'hA0;
mem[16'h0A09] = 8'hA0;
mem[16'h0A0A] = 8'hA0;
mem[16'h0A0B] = 8'hA0;
mem[16'h0A0C] = 8'hA0;
mem[16'h0A0D] = 8'hA0;
mem[16'h0A0E] = 8'hA0;
mem[16'h0A0F] = 8'hA0;
mem[16'h0A10] = 8'hA0;
mem[16'h0A11] = 8'hA0;
mem[16'h0A12] = 8'hA0;
mem[16'h0A13] = 8'hA0;
mem[16'h0A14] = 8'hA0;
mem[16'h0A15] = 8'hA0;
mem[16'h0A16] = 8'hA0;
mem[16'h0A17] = 8'hA0;
mem[16'h0A18] = 8'hA0;
mem[16'h0A19] = 8'hA0;
mem[16'h0A1A] = 8'hA0;
mem[16'h0A1B] = 8'hA0;
mem[16'h0A1C] = 8'hA0;
mem[16'h0A1D] = 8'hA0;
mem[16'h0A1E] = 8'hA0;
mem[16'h0A1F] = 8'hA0;
mem[16'h0A20] = 8'hA0;
mem[16'h0A21] = 8'hA0;
mem[16'h0A22] = 8'hA0;
mem[16'h0A23] = 8'hA0;
mem[16'h0A24] = 8'hA0;
mem[16'h0A25] = 8'hAA;
mem[16'h0A26] = 8'hAA;
mem[16'h0A27] = 8'hA0;
mem[16'h0A28] = 8'hAA;
mem[16'h0A29] = 8'hAA;
mem[16'h0A2A] = 8'hA0;
mem[16'h0A2B] = 8'hA0;
mem[16'h0A2C] = 8'hA0;
mem[16'h0A2D] = 8'hA0;
mem[16'h0A2E] = 8'hA0;
mem[16'h0A2F] = 8'hA0;
mem[16'h0A30] = 8'hA0;
mem[16'h0A31] = 8'hA0;
mem[16'h0A32] = 8'hA0;
mem[16'h0A33] = 8'hA0;
mem[16'h0A34] = 8'hA0;
mem[16'h0A35] = 8'hA0;
mem[16'h0A36] = 8'hA0;
mem[16'h0A37] = 8'hA0;
mem[16'h0A38] = 8'hA0;
mem[16'h0A39] = 8'hA0;
mem[16'h0A3A] = 8'hA0;
mem[16'h0A3B] = 8'hA0;
mem[16'h0A3C] = 8'hA0;
mem[16'h0A3D] = 8'hA0;
mem[16'h0A3E] = 8'hA0;
mem[16'h0A3F] = 8'hA0;
mem[16'h0A40] = 8'hA0;
mem[16'h0A41] = 8'hA0;
mem[16'h0A42] = 8'hA0;
mem[16'h0A43] = 8'hA0;
mem[16'h0A44] = 8'hA0;
mem[16'h0A45] = 8'hA0;
mem[16'h0A46] = 8'hA0;
mem[16'h0A47] = 8'hA0;
mem[16'h0A48] = 8'hA0;
mem[16'h0A49] = 8'hA0;
mem[16'h0A4A] = 8'hA0;
mem[16'h0A4B] = 8'hA0;
mem[16'h0A4C] = 8'hA0;
mem[16'h0A4D] = 8'hAA;
mem[16'h0A4E] = 8'hAA;
mem[16'h0A4F] = 8'hA0;
mem[16'h0A50] = 8'hAA;
mem[16'h0A51] = 8'hAA;
mem[16'h0A52] = 8'hA0;
mem[16'h0A53] = 8'hA0;
mem[16'h0A54] = 8'hA0;
mem[16'h0A55] = 8'hA0;
mem[16'h0A56] = 8'hA0;
mem[16'h0A57] = 8'hA0;
mem[16'h0A58] = 8'hA0;
mem[16'h0A59] = 8'hA0;
mem[16'h0A5A] = 8'hA0;
mem[16'h0A5B] = 8'hA0;
mem[16'h0A5C] = 8'hA0;
mem[16'h0A5D] = 8'hA0;
mem[16'h0A5E] = 8'hA0;
mem[16'h0A5F] = 8'hA0;
mem[16'h0A60] = 8'hA0;
mem[16'h0A61] = 8'hA0;
mem[16'h0A62] = 8'hA0;
mem[16'h0A63] = 8'hA0;
mem[16'h0A64] = 8'hA0;
mem[16'h0A65] = 8'hA0;
mem[16'h0A66] = 8'hA0;
mem[16'h0A67] = 8'hA0;
mem[16'h0A68] = 8'hA0;
mem[16'h0A69] = 8'hA0;
mem[16'h0A6A] = 8'hA0;
mem[16'h0A6B] = 8'hA0;
mem[16'h0A6C] = 8'hA0;
mem[16'h0A6D] = 8'hA0;
mem[16'h0A6E] = 8'hA0;
mem[16'h0A6F] = 8'hA0;
mem[16'h0A70] = 8'hA0;
mem[16'h0A71] = 8'hA0;
mem[16'h0A72] = 8'hA0;
mem[16'h0A73] = 8'hA0;
mem[16'h0A74] = 8'hA0;
mem[16'h0A75] = 8'hAA;
mem[16'h0A76] = 8'hAA;
mem[16'h0A77] = 8'hA0;
mem[16'h0A78] = 8'h60;
mem[16'h0A79] = 8'h42;
mem[16'h0A7A] = 8'h42;
mem[16'h0A7B] = 8'h42;
mem[16'h0A7C] = 8'h42;
mem[16'h0A7D] = 8'h42;
mem[16'h0A7E] = 8'h3C;
mem[16'h0A7F] = 8'h00;
mem[16'h0A80] = 8'hAA;
mem[16'h0A81] = 8'hAA;
mem[16'h0A82] = 8'hA0;
mem[16'h0A83] = 8'hA0;
mem[16'h0A84] = 8'hA0;
mem[16'h0A85] = 8'hA0;
mem[16'h0A86] = 8'hA0;
mem[16'h0A87] = 8'hA0;
mem[16'h0A88] = 8'hA0;
mem[16'h0A89] = 8'hA0;
mem[16'h0A8A] = 8'hA0;
mem[16'h0A8B] = 8'hC2;
mem[16'h0A8C] = 8'hD9;
mem[16'h0A8D] = 8'hA0;
mem[16'h0A8E] = 8'hCF;
mem[16'h0A8F] = 8'hCC;
mem[16'h0A90] = 8'hC1;
mem[16'h0A91] = 8'hC6;
mem[16'h0A92] = 8'hA0;
mem[16'h0A93] = 8'hCC;
mem[16'h0A94] = 8'hD5;
mem[16'h0A95] = 8'hC2;
mem[16'h0A96] = 8'hC5;
mem[16'h0A97] = 8'hC3;
mem[16'h0A98] = 8'hCB;
mem[16'h0A99] = 8'hA0;
mem[16'h0A9A] = 8'hA0;
mem[16'h0A9B] = 8'hA0;
mem[16'h0A9C] = 8'hA0;
mem[16'h0A9D] = 8'hA0;
mem[16'h0A9E] = 8'hA0;
mem[16'h0A9F] = 8'hA0;
mem[16'h0AA0] = 8'hA0;
mem[16'h0AA1] = 8'hA0;
mem[16'h0AA2] = 8'hA0;
mem[16'h0AA3] = 8'hA0;
mem[16'h0AA4] = 8'hA0;
mem[16'h0AA5] = 8'hAA;
mem[16'h0AA6] = 8'hAA;
mem[16'h0AA7] = 8'hA0;
mem[16'h0AA8] = 8'hAA;
mem[16'h0AA9] = 8'hAA;
mem[16'h0AAA] = 8'hA0;
mem[16'h0AAB] = 8'hA0;
mem[16'h0AAC] = 8'h13;
mem[16'h0AAD] = 8'h10;
mem[16'h0AAE] = 8'h01;
mem[16'h0AAF] = 8'h03;
mem[16'h0AB0] = 8'h05;
mem[16'h0AB1] = 8'h20;
mem[16'h0AB2] = 8'h02;
mem[16'h0AB3] = 8'h01;
mem[16'h0AB4] = 8'h12;
mem[16'h0AB5] = 8'hA0;
mem[16'h0AB6] = 8'hD4;
mem[16'h0AB7] = 8'hCF;
mem[16'h0AB8] = 8'hA0;
mem[16'h0AB9] = 8'hD3;
mem[16'h0ABA] = 8'hD4;
mem[16'h0ABB] = 8'hC1;
mem[16'h0ABC] = 8'hD2;
mem[16'h0ABD] = 8'hD4;
mem[16'h0ABE] = 8'hA0;
mem[16'h0ABF] = 8'hC6;
mem[16'h0AC0] = 8'hD2;
mem[16'h0AC1] = 8'hCF;
mem[16'h0AC2] = 8'hC7;
mem[16'h0AC3] = 8'hC7;
mem[16'h0AC4] = 8'hC9;
mem[16'h0AC5] = 8'hCE;
mem[16'h0AC6] = 8'hC7;
mem[16'h0AC7] = 8'hA0;
mem[16'h0AC8] = 8'hA0;
mem[16'h0AC9] = 8'hA0;
mem[16'h0ACA] = 8'hA0;
mem[16'h0ACB] = 8'hA0;
mem[16'h0ACC] = 8'hA0;
mem[16'h0ACD] = 8'hAA;
mem[16'h0ACE] = 8'hAA;
mem[16'h0ACF] = 8'hA0;
mem[16'h0AD0] = 8'hAA;
mem[16'h0AD1] = 8'hAA;
mem[16'h0AD2] = 8'hAA;
mem[16'h0AD3] = 8'hAA;
mem[16'h0AD4] = 8'hAA;
mem[16'h0AD5] = 8'hAA;
mem[16'h0AD6] = 8'hAA;
mem[16'h0AD7] = 8'hAA;
mem[16'h0AD8] = 8'hAA;
mem[16'h0AD9] = 8'hAA;
mem[16'h0ADA] = 8'hAA;
mem[16'h0ADB] = 8'hAA;
mem[16'h0ADC] = 8'hAA;
mem[16'h0ADD] = 8'hAA;
mem[16'h0ADE] = 8'hAA;
mem[16'h0ADF] = 8'hAA;
mem[16'h0AE0] = 8'hAA;
mem[16'h0AE1] = 8'hAA;
mem[16'h0AE2] = 8'hAA;
mem[16'h0AE3] = 8'hAA;
mem[16'h0AE4] = 8'hAA;
mem[16'h0AE5] = 8'hAA;
mem[16'h0AE6] = 8'hAA;
mem[16'h0AE7] = 8'hAA;
mem[16'h0AE8] = 8'hAA;
mem[16'h0AE9] = 8'hAA;
mem[16'h0AEA] = 8'hAA;
mem[16'h0AEB] = 8'hAA;
mem[16'h0AEC] = 8'hAA;
mem[16'h0AED] = 8'hAA;
mem[16'h0AEE] = 8'hAA;
mem[16'h0AEF] = 8'hAA;
mem[16'h0AF0] = 8'hAA;
mem[16'h0AF1] = 8'hAA;
mem[16'h0AF2] = 8'hAA;
mem[16'h0AF3] = 8'hAA;
mem[16'h0AF4] = 8'hAA;
mem[16'h0AF5] = 8'hAA;
mem[16'h0AF6] = 8'hAA;
mem[16'h0AF7] = 8'hA0;
mem[16'h0AF8] = 8'h02;
mem[16'h0AF9] = 8'h00;
mem[16'h0AFA] = 8'h00;
mem[16'h0AFB] = 8'h00;
mem[16'h0AFC] = 8'h00;
mem[16'h0AFD] = 8'h00;
mem[16'h0AFE] = 8'h00;
mem[16'h0AFF] = 8'hFF;
mem[16'h0B00] = 8'hAA;
mem[16'h0B01] = 8'hAA;
mem[16'h0B02] = 8'hA0;
mem[16'h0B03] = 8'hA0;
mem[16'h0B04] = 8'hA0;
mem[16'h0B05] = 8'hA0;
mem[16'h0B06] = 8'hA0;
mem[16'h0B07] = 8'hA0;
mem[16'h0B08] = 8'hA0;
mem[16'h0B09] = 8'hA0;
mem[16'h0B0A] = 8'hA0;
mem[16'h0B0B] = 8'hA0;
mem[16'h0B0C] = 8'hA0;
mem[16'h0B0D] = 8'hA0;
mem[16'h0B0E] = 8'hA0;
mem[16'h0B0F] = 8'hA0;
mem[16'h0B10] = 8'hA0;
mem[16'h0B11] = 8'hA0;
mem[16'h0B12] = 8'hA0;
mem[16'h0B13] = 8'hA0;
mem[16'h0B14] = 8'hA0;
mem[16'h0B15] = 8'hA0;
mem[16'h0B16] = 8'hA0;
mem[16'h0B17] = 8'hA0;
mem[16'h0B18] = 8'hA0;
mem[16'h0B19] = 8'hA0;
mem[16'h0B1A] = 8'hA0;
mem[16'h0B1B] = 8'hA0;
mem[16'h0B1C] = 8'hA0;
mem[16'h0B1D] = 8'hA0;
mem[16'h0B1E] = 8'hA0;
mem[16'h0B1F] = 8'hA0;
mem[16'h0B20] = 8'hA0;
mem[16'h0B21] = 8'hA0;
mem[16'h0B22] = 8'hA0;
mem[16'h0B23] = 8'hA0;
mem[16'h0B24] = 8'hA0;
mem[16'h0B25] = 8'hAA;
mem[16'h0B26] = 8'hAA;
mem[16'h0B27] = 8'hA0;
mem[16'h0B28] = 8'hAA;
mem[16'h0B29] = 8'hAA;
mem[16'h0B2A] = 8'hA0;
mem[16'h0B2B] = 8'hA0;
mem[16'h0B2C] = 8'hA0;
mem[16'h0B2D] = 8'hA0;
mem[16'h0B2E] = 8'hA0;
mem[16'h0B2F] = 8'hA0;
mem[16'h0B30] = 8'hA0;
mem[16'h0B31] = 8'hA0;
mem[16'h0B32] = 8'hA0;
mem[16'h0B33] = 8'hA0;
mem[16'h0B34] = 8'hA0;
mem[16'h0B35] = 8'hA0;
mem[16'h0B36] = 8'hA0;
mem[16'h0B37] = 8'hA0;
mem[16'h0B38] = 8'hA0;
mem[16'h0B39] = 8'hA0;
mem[16'h0B3A] = 8'hA0;
mem[16'h0B3B] = 8'hA0;
mem[16'h0B3C] = 8'hA0;
mem[16'h0B3D] = 8'hA0;
mem[16'h0B3E] = 8'hA0;
mem[16'h0B3F] = 8'hA0;
mem[16'h0B40] = 8'hA0;
mem[16'h0B41] = 8'hA0;
mem[16'h0B42] = 8'hA0;
mem[16'h0B43] = 8'hA0;
mem[16'h0B44] = 8'hA0;
mem[16'h0B45] = 8'hA0;
mem[16'h0B46] = 8'hA0;
mem[16'h0B47] = 8'hA0;
mem[16'h0B48] = 8'hA0;
mem[16'h0B49] = 8'hA0;
mem[16'h0B4A] = 8'hA0;
mem[16'h0B4B] = 8'hA0;
mem[16'h0B4C] = 8'hA0;
mem[16'h0B4D] = 8'hAA;
mem[16'h0B4E] = 8'hAA;
mem[16'h0B4F] = 8'hA0;
mem[16'h0B50] = 8'hA0;
mem[16'h0B51] = 8'hA0;
mem[16'h0B52] = 8'hA0;
mem[16'h0B53] = 8'hA0;
mem[16'h0B54] = 8'hA0;
mem[16'h0B55] = 8'hA0;
mem[16'h0B56] = 8'hA0;
mem[16'h0B57] = 8'hA0;
mem[16'h0B58] = 8'hA0;
mem[16'h0B59] = 8'hA0;
mem[16'h0B5A] = 8'hA0;
mem[16'h0B5B] = 8'hA0;
mem[16'h0B5C] = 8'hA0;
mem[16'h0B5D] = 8'hA0;
mem[16'h0B5E] = 8'hA0;
mem[16'h0B5F] = 8'hA0;
mem[16'h0B60] = 8'hA0;
mem[16'h0B61] = 8'hA0;
mem[16'h0B62] = 8'hA0;
mem[16'h0B63] = 8'hA0;
mem[16'h0B64] = 8'hA0;
mem[16'h0B65] = 8'hA0;
mem[16'h0B66] = 8'hA0;
mem[16'h0B67] = 8'hA0;
mem[16'h0B68] = 8'hA0;
mem[16'h0B69] = 8'hA0;
mem[16'h0B6A] = 8'hA0;
mem[16'h0B6B] = 8'hA0;
mem[16'h0B6C] = 8'hA0;
mem[16'h0B6D] = 8'hA0;
mem[16'h0B6E] = 8'hA0;
mem[16'h0B6F] = 8'hA0;
mem[16'h0B70] = 8'hA0;
mem[16'h0B71] = 8'hA0;
mem[16'h0B72] = 8'hA0;
mem[16'h0B73] = 8'hA0;
mem[16'h0B74] = 8'hA0;
mem[16'h0B75] = 8'hA0;
mem[16'h0B76] = 8'hA0;
mem[16'h0B77] = 8'hA0;
mem[16'h0B78] = 8'h00;
mem[16'h0B79] = 8'h00;
mem[16'h0B7A] = 8'h38;
mem[16'h0B7B] = 8'h44;
mem[16'h0B7C] = 8'h44;
mem[16'h0B7D] = 8'h44;
mem[16'h0B7E] = 8'h38;
mem[16'h0B7F] = 8'h00;
mem[16'h0B80] = 8'hAA;
mem[16'h0B81] = 8'hAA;
mem[16'h0B82] = 8'hA0;
mem[16'h0B83] = 8'hA0;
mem[16'h0B84] = 8'hA0;
mem[16'h0B85] = 8'hA0;
mem[16'h0B86] = 8'hA0;
mem[16'h0B87] = 8'hA0;
mem[16'h0B88] = 8'hCD;
mem[16'h0B89] = 8'hC1;
mem[16'h0B8A] = 8'hC9;
mem[16'h0B8B] = 8'hCE;
mem[16'h0B8C] = 8'hA0;
mem[16'h0B8D] = 8'hD3;
mem[16'h0B8E] = 8'hD4;
mem[16'h0B8F] = 8'hD2;
mem[16'h0B90] = 8'hC5;
mem[16'h0B91] = 8'hC5;
mem[16'h0B92] = 8'hD4;
mem[16'h0B93] = 8'hA0;
mem[16'h0B94] = 8'hD0;
mem[16'h0B95] = 8'hD5;
mem[16'h0B96] = 8'hC2;
mem[16'h0B97] = 8'hCC;
mem[16'h0B98] = 8'hC9;
mem[16'h0B99] = 8'hD3;
mem[16'h0B9A] = 8'hC8;
mem[16'h0B9B] = 8'hC9;
mem[16'h0B9C] = 8'hCE;
mem[16'h0B9D] = 8'hC7;
mem[16'h0B9E] = 8'hA0;
mem[16'h0B9F] = 8'hA0;
mem[16'h0BA0] = 8'hA0;
mem[16'h0BA1] = 8'hA0;
mem[16'h0BA2] = 8'hA0;
mem[16'h0BA3] = 8'hA0;
mem[16'h0BA4] = 8'hA0;
mem[16'h0BA5] = 8'hAA;
mem[16'h0BA6] = 8'hAA;
mem[16'h0BA7] = 8'hA0;
mem[16'h0BA8] = 8'hAA;
mem[16'h0BA9] = 8'hAA;
mem[16'h0BAA] = 8'hA0;
mem[16'h0BAB] = 8'hA0;
mem[16'h0BAC] = 8'h04;
mem[16'h0BAD] = 8'hA0;
mem[16'h0BAE] = 8'hD4;
mem[16'h0BAF] = 8'hCF;
mem[16'h0BB0] = 8'hA0;
mem[16'h0BB1] = 8'hC4;
mem[16'h0BB2] = 8'hC5;
mem[16'h0BB3] = 8'hC6;
mem[16'h0BB4] = 8'hC9;
mem[16'h0BB5] = 8'hCE;
mem[16'h0BB6] = 8'hC5;
mem[16'h0BB7] = 8'hA0;
mem[16'h0BB8] = 8'hD9;
mem[16'h0BB9] = 8'hCF;
mem[16'h0BBA] = 8'hD5;
mem[16'h0BBB] = 8'hD2;
mem[16'h0BBC] = 8'hA0;
mem[16'h0BBD] = 8'hCF;
mem[16'h0BBE] = 8'hD7;
mem[16'h0BBF] = 8'hCE;
mem[16'h0BC0] = 8'hA0;
mem[16'h0BC1] = 8'hCB;
mem[16'h0BC2] = 8'hC5;
mem[16'h0BC3] = 8'hD9;
mem[16'h0BC4] = 8'hD3;
mem[16'h0BC5] = 8'hA0;
mem[16'h0BC6] = 8'hA0;
mem[16'h0BC7] = 8'hA0;
mem[16'h0BC8] = 8'hA0;
mem[16'h0BC9] = 8'hA0;
mem[16'h0BCA] = 8'hA0;
mem[16'h0BCB] = 8'hA0;
mem[16'h0BCC] = 8'hA0;
mem[16'h0BCD] = 8'hAA;
mem[16'h0BCE] = 8'hAA;
mem[16'h0BCF] = 8'hA0;
mem[16'h0BD0] = 8'hA0;
mem[16'h0BD1] = 8'hA0;
mem[16'h0BD2] = 8'hA0;
mem[16'h0BD3] = 8'hA0;
mem[16'h0BD4] = 8'hA0;
mem[16'h0BD5] = 8'hA0;
mem[16'h0BD6] = 8'hA0;
mem[16'h0BD7] = 8'hA0;
mem[16'h0BD8] = 8'hA0;
mem[16'h0BD9] = 8'hA0;
mem[16'h0BDA] = 8'hA0;
mem[16'h0BDB] = 8'hA0;
mem[16'h0BDC] = 8'hA0;
mem[16'h0BDD] = 8'hA0;
mem[16'h0BDE] = 8'hA0;
mem[16'h0BDF] = 8'hA0;
mem[16'h0BE0] = 8'hA0;
mem[16'h0BE1] = 8'hA0;
mem[16'h0BE2] = 8'hA0;
mem[16'h0BE3] = 8'hA0;
mem[16'h0BE4] = 8'hA0;
mem[16'h0BE5] = 8'hA0;
mem[16'h0BE6] = 8'hA0;
mem[16'h0BE7] = 8'hA0;
mem[16'h0BE8] = 8'hA0;
mem[16'h0BE9] = 8'hA0;
mem[16'h0BEA] = 8'hA0;
mem[16'h0BEB] = 8'hA0;
mem[16'h0BEC] = 8'hA0;
mem[16'h0BED] = 8'hA0;
mem[16'h0BEE] = 8'hA0;
mem[16'h0BEF] = 8'hA0;
mem[16'h0BF0] = 8'hA0;
mem[16'h0BF1] = 8'hA0;
mem[16'h0BF2] = 8'hA0;
mem[16'h0BF3] = 8'hA0;
mem[16'h0BF4] = 8'hA0;
mem[16'h0BF5] = 8'hA0;
mem[16'h0BF6] = 8'hA0;
mem[16'h0BF7] = 8'hA0;
mem[16'h0BF8] = 8'hFF;
mem[16'h0BF9] = 8'hFF;
mem[16'h0BFA] = 8'hFF;
mem[16'h0BFB] = 8'hFF;
mem[16'h0BFC] = 8'hFF;
mem[16'h0BFD] = 8'h0F;
mem[16'h0BFE] = 8'hAB;
mem[16'h0BFF] = 8'hDC;
mem[16'h0C00] = 8'hA9;
mem[16'h0C01] = 8'h00;
mem[16'h0C02] = 8'h85;
mem[16'h0C03] = 8'h00;
mem[16'h0C04] = 8'h85;
mem[16'h0C05] = 8'h02;
mem[16'h0C06] = 8'hA9;
mem[16'h0C07] = 8'h16;
mem[16'h0C08] = 8'h85;
mem[16'h0C09] = 8'h01;
mem[16'h0C0A] = 8'hA9;
mem[16'h0C0B] = 8'h96;
mem[16'h0C0C] = 8'h85;
mem[16'h0C0D] = 8'h03;
mem[16'h0C0E] = 8'hA0;
mem[16'h0C0F] = 8'h00;
mem[16'h0C10] = 8'hB1;
mem[16'h0C11] = 8'h00;
mem[16'h0C12] = 8'h91;
mem[16'h0C13] = 8'h02;
mem[16'h0C14] = 8'hC8;
mem[16'h0C15] = 8'hD0;
mem[16'h0C16] = 8'hF9;
mem[16'h0C17] = 8'hE6;
mem[16'h0C18] = 8'h01;
mem[16'h0C19] = 8'hE6;
mem[16'h0C1A] = 8'h03;
mem[16'h0C1B] = 8'hA5;
mem[16'h0C1C] = 8'h03;
mem[16'h0C1D] = 8'hC9;
mem[16'h0C1E] = 8'hC0;
mem[16'h0C1F] = 8'hD0;
mem[16'h0C20] = 8'hEF;
mem[16'h0C21] = 8'hEA;
mem[16'h0C22] = 8'hA2;
mem[16'h0C23] = 8'h00;
mem[16'h0C24] = 8'hBD;
mem[16'h0C25] = 8'h00;
mem[16'h0C26] = 8'h0E;
mem[16'h0C27] = 8'h95;
mem[16'h0C28] = 8'h00;
mem[16'h0C29] = 8'hBD;
mem[16'h0C2A] = 8'h00;
mem[16'h0C2B] = 8'h0F;
mem[16'h0C2C] = 8'h9D;
mem[16'h0C2D] = 8'h00;
mem[16'h0C2E] = 8'h01;
mem[16'h0C2F] = 8'hBD;
mem[16'h0C30] = 8'h00;
mem[16'h0C31] = 8'h10;
mem[16'h0C32] = 8'h9D;
mem[16'h0C33] = 8'h00;
mem[16'h0C34] = 8'h02;
mem[16'h0C35] = 8'hBD;
mem[16'h0C36] = 8'h00;
mem[16'h0C37] = 8'h11;
mem[16'h0C38] = 8'h9D;
mem[16'h0C39] = 8'h00;
mem[16'h0C3A] = 8'h03;
mem[16'h0C3B] = 8'hBD;
mem[16'h0C3C] = 8'h00;
mem[16'h0C3D] = 8'h12;
mem[16'h0C3E] = 8'h9D;
mem[16'h0C3F] = 8'h00;
mem[16'h0C40] = 8'h04;
mem[16'h0C41] = 8'hBD;
mem[16'h0C42] = 8'h00;
mem[16'h0C43] = 8'h13;
mem[16'h0C44] = 8'h9D;
mem[16'h0C45] = 8'h00;
mem[16'h0C46] = 8'h05;
mem[16'h0C47] = 8'hBD;
mem[16'h0C48] = 8'h00;
mem[16'h0C49] = 8'h14;
mem[16'h0C4A] = 8'h9D;
mem[16'h0C4B] = 8'h00;
mem[16'h0C4C] = 8'h06;
mem[16'h0C4D] = 8'hBD;
mem[16'h0C4E] = 8'h00;
mem[16'h0C4F] = 8'h15;
mem[16'h0C50] = 8'h9D;
mem[16'h0C51] = 8'h00;
mem[16'h0C52] = 8'h07;
mem[16'h0C53] = 8'hE8;
mem[16'h0C54] = 8'hD0;
mem[16'h0C55] = 8'hCE;
mem[16'h0C56] = 8'hEA;
mem[16'h0C57] = 8'h4C;
mem[16'h0C58] = 8'h00;
mem[16'h0C59] = 8'h9C;
mem[16'h0C5A] = 8'hC9;
mem[16'h0C5B] = 8'hD8;
mem[16'h0C5C] = 8'hD0;
mem[16'h0C5D] = 8'h32;
mem[16'h0C5E] = 8'hAD;
mem[16'h0C5F] = 8'h98;
mem[16'h0C60] = 8'h0B;
mem[16'h0C61] = 8'hC9;
mem[16'h0C62] = 8'hC5;
mem[16'h0C63] = 8'hD0;
mem[16'h0C64] = 8'h2B;
mem[16'h0C65] = 8'hAD;
mem[16'h0C66] = 8'h99;
mem[16'h0C67] = 8'h0B;
mem[16'h0C68] = 8'hC9;
mem[16'h0C69] = 8'hD2;
mem[16'h0C6A] = 8'hD0;
mem[16'h0C6B] = 8'h24;
mem[16'h0C6C] = 8'hAD;
mem[16'h0C6D] = 8'h9A;
mem[16'h0C6E] = 8'h0B;
mem[16'h0C6F] = 8'hC9;
mem[16'h0C70] = 8'hCF;
mem[16'h0C71] = 8'hD0;
mem[16'h0C72] = 8'h1D;
mem[16'h0C73] = 8'hAD;
mem[16'h0C74] = 8'h9B;
mem[16'h0C75] = 8'h0B;
mem[16'h0C76] = 8'hC9;
mem[16'h0C77] = 8'hD8;
mem[16'h0C78] = 8'hD0;
mem[16'h0C79] = 8'h16;
mem[16'h0C7A] = 8'h4C;
mem[16'h0C7B] = 8'h00;
mem[16'h0C7C] = 8'h9C;
mem[16'h0C7D] = 8'hDC;
mem[16'h0C7E] = 8'hDC;
mem[16'h0C7F] = 8'hDC;
mem[16'h0C80] = 8'hDC;
mem[16'h0C81] = 8'hDC;
mem[16'h0C82] = 8'hDC;
mem[16'h0C83] = 8'hDC;
mem[16'h0C84] = 8'hDC;
mem[16'h0C85] = 8'hDC;
mem[16'h0C86] = 8'hDC;
mem[16'h0C87] = 8'hDC;
mem[16'h0C88] = 8'hDC;
mem[16'h0C89] = 8'hDC;
mem[16'h0C8A] = 8'hDC;
mem[16'h0C8B] = 8'hDC;
mem[16'h0C8C] = 8'hDC;
mem[16'h0C8D] = 8'hDC;
mem[16'h0C8E] = 8'hDC;
mem[16'h0C8F] = 8'hDC;
mem[16'h0C90] = 8'h4C;
mem[16'h0C91] = 8'h00;
mem[16'h0C92] = 8'hC6;
mem[16'h0C93] = 8'hDC;
mem[16'h0C94] = 8'hDC;
mem[16'h0C95] = 8'hDC;
mem[16'h0C96] = 8'hDC;
mem[16'h0C97] = 8'hDC;
mem[16'h0C98] = 8'hDC;
mem[16'h0C99] = 8'hDC;
mem[16'h0C9A] = 8'hDC;
mem[16'h0C9B] = 8'hDC;
mem[16'h0C9C] = 8'hDC;
mem[16'h0C9D] = 8'hDC;
mem[16'h0C9E] = 8'hDC;
mem[16'h0C9F] = 8'hDC;
mem[16'h0CA0] = 8'hDC;
mem[16'h0CA1] = 8'hDC;
mem[16'h0CA2] = 8'hDC;
mem[16'h0CA3] = 8'hDC;
mem[16'h0CA4] = 8'hDC;
mem[16'h0CA5] = 8'hDC;
mem[16'h0CA6] = 8'hDC;
mem[16'h0CA7] = 8'hDC;
mem[16'h0CA8] = 8'hDC;
mem[16'h0CA9] = 8'hDC;
mem[16'h0CAA] = 8'hDC;
mem[16'h0CAB] = 8'hDC;
mem[16'h0CAC] = 8'hDC;
mem[16'h0CAD] = 8'hDC;
mem[16'h0CAE] = 8'hDC;
mem[16'h0CAF] = 8'hDC;
mem[16'h0CB0] = 8'hDC;
mem[16'h0CB1] = 8'hDC;
mem[16'h0CB2] = 8'hDC;
mem[16'h0CB3] = 8'hDC;
mem[16'h0CB4] = 8'hDC;
mem[16'h0CB5] = 8'hDC;
mem[16'h0CB6] = 8'hDC;
mem[16'h0CB7] = 8'hDC;
mem[16'h0CB8] = 8'hDC;
mem[16'h0CB9] = 8'hDC;
mem[16'h0CBA] = 8'hDC;
mem[16'h0CBB] = 8'hDC;
mem[16'h0CBC] = 8'hDC;
mem[16'h0CBD] = 8'hDC;
mem[16'h0CBE] = 8'hDC;
mem[16'h0CBF] = 8'hDC;
mem[16'h0CC0] = 8'hDC;
mem[16'h0CC1] = 8'hDC;
mem[16'h0CC2] = 8'hDC;
mem[16'h0CC3] = 8'hDC;
mem[16'h0CC4] = 8'hDC;
mem[16'h0CC5] = 8'hDC;
mem[16'h0CC6] = 8'hDC;
mem[16'h0CC7] = 8'hDC;
mem[16'h0CC8] = 8'hDC;
mem[16'h0CC9] = 8'hDC;
mem[16'h0CCA] = 8'hDC;
mem[16'h0CCB] = 8'hDC;
mem[16'h0CCC] = 8'hDC;
mem[16'h0CCD] = 8'hDC;
mem[16'h0CCE] = 8'hDC;
mem[16'h0CCF] = 8'hDC;
mem[16'h0CD0] = 8'hDC;
mem[16'h0CD1] = 8'hDC;
mem[16'h0CD2] = 8'hDC;
mem[16'h0CD3] = 8'hDC;
mem[16'h0CD4] = 8'hDC;
mem[16'h0CD5] = 8'hDC;
mem[16'h0CD6] = 8'hDC;
mem[16'h0CD7] = 8'hDC;
mem[16'h0CD8] = 8'hDC;
mem[16'h0CD9] = 8'hDC;
mem[16'h0CDA] = 8'hDC;
mem[16'h0CDB] = 8'hDC;
mem[16'h0CDC] = 8'hDC;
mem[16'h0CDD] = 8'hDC;
mem[16'h0CDE] = 8'hDC;
mem[16'h0CDF] = 8'hDC;
mem[16'h0CE0] = 8'hDC;
mem[16'h0CE1] = 8'hDC;
mem[16'h0CE2] = 8'hDC;
mem[16'h0CE3] = 8'hDC;
mem[16'h0CE4] = 8'hDC;
mem[16'h0CE5] = 8'hDC;
mem[16'h0CE6] = 8'hDC;
mem[16'h0CE7] = 8'hDC;
mem[16'h0CE8] = 8'hDC;
mem[16'h0CE9] = 8'hDC;
mem[16'h0CEA] = 8'hDC;
mem[16'h0CEB] = 8'hDC;
mem[16'h0CEC] = 8'hDC;
mem[16'h0CED] = 8'hDC;
mem[16'h0CEE] = 8'hDC;
mem[16'h0CEF] = 8'hDC;
mem[16'h0CF0] = 8'hDC;
mem[16'h0CF1] = 8'hDC;
mem[16'h0CF2] = 8'hDC;
mem[16'h0CF3] = 8'hDC;
mem[16'h0CF4] = 8'hDC;
mem[16'h0CF5] = 8'hDC;
mem[16'h0CF6] = 8'hDC;
mem[16'h0CF7] = 8'hDC;
mem[16'h0CF8] = 8'hDC;
mem[16'h0CF9] = 8'hDC;
mem[16'h0CFA] = 8'hDC;
mem[16'h0CFB] = 8'hDC;
mem[16'h0CFC] = 8'hDC;
mem[16'h0CFD] = 8'hDC;
mem[16'h0CFE] = 8'hDC;
mem[16'h0CFF] = 8'hDC;
mem[16'h0D00] = 8'hAD;
mem[16'h0D01] = 8'h55;
mem[16'h0D02] = 8'hC0;
mem[16'h0D03] = 8'hAD;
mem[16'h0D04] = 8'h52;
mem[16'h0D05] = 8'hC0;
mem[16'h0D06] = 8'hAD;
mem[16'h0D07] = 8'h51;
mem[16'h0D08] = 8'hC0;
mem[16'h0D09] = 8'h60;
mem[16'h0D0A] = 8'hDC;
mem[16'h0D0B] = 8'hDC;
mem[16'h0D0C] = 8'hDC;
mem[16'h0D0D] = 8'hDC;
mem[16'h0D0E] = 8'hDC;
mem[16'h0D0F] = 8'hDC;
mem[16'h0D10] = 8'hDC;
mem[16'h0D11] = 8'hDC;
mem[16'h0D12] = 8'hDC;
mem[16'h0D13] = 8'hDC;
mem[16'h0D14] = 8'hDC;
mem[16'h0D15] = 8'hDC;
mem[16'h0D16] = 8'hDC;
mem[16'h0D17] = 8'hDC;
mem[16'h0D18] = 8'hDC;
mem[16'h0D19] = 8'hDC;
mem[16'h0D1A] = 8'hDC;
mem[16'h0D1B] = 8'hDC;
mem[16'h0D1C] = 8'hDC;
mem[16'h0D1D] = 8'hDC;
mem[16'h0D1E] = 8'hDC;
mem[16'h0D1F] = 8'hDC;
mem[16'h0D20] = 8'hDC;
mem[16'h0D21] = 8'hDC;
mem[16'h0D22] = 8'hDC;
mem[16'h0D23] = 8'hDC;
mem[16'h0D24] = 8'hDC;
mem[16'h0D25] = 8'hDC;
mem[16'h0D26] = 8'hDC;
mem[16'h0D27] = 8'hDC;
mem[16'h0D28] = 8'hDC;
mem[16'h0D29] = 8'hDC;
mem[16'h0D2A] = 8'hDC;
mem[16'h0D2B] = 8'hDC;
mem[16'h0D2C] = 8'hDC;
mem[16'h0D2D] = 8'hDC;
mem[16'h0D2E] = 8'hDC;
mem[16'h0D2F] = 8'hDC;
mem[16'h0D30] = 8'hDC;
mem[16'h0D31] = 8'hDC;
mem[16'h0D32] = 8'hDC;
mem[16'h0D33] = 8'hDC;
mem[16'h0D34] = 8'hDC;
mem[16'h0D35] = 8'hDC;
mem[16'h0D36] = 8'hDC;
mem[16'h0D37] = 8'hDC;
mem[16'h0D38] = 8'hDC;
mem[16'h0D39] = 8'hDC;
mem[16'h0D3A] = 8'hDC;
mem[16'h0D3B] = 8'hDC;
mem[16'h0D3C] = 8'hDC;
mem[16'h0D3D] = 8'hDC;
mem[16'h0D3E] = 8'hDC;
mem[16'h0D3F] = 8'hDC;
mem[16'h0D40] = 8'hDC;
mem[16'h0D41] = 8'hDC;
mem[16'h0D42] = 8'hDC;
mem[16'h0D43] = 8'hDC;
mem[16'h0D44] = 8'hDC;
mem[16'h0D45] = 8'hDC;
mem[16'h0D46] = 8'hDC;
mem[16'h0D47] = 8'hDC;
mem[16'h0D48] = 8'hDC;
mem[16'h0D49] = 8'hDC;
mem[16'h0D4A] = 8'hDC;
mem[16'h0D4B] = 8'hDC;
mem[16'h0D4C] = 8'hDC;
mem[16'h0D4D] = 8'hDC;
mem[16'h0D4E] = 8'hDC;
mem[16'h0D4F] = 8'hDC;
mem[16'h0D50] = 8'hDC;
mem[16'h0D51] = 8'hDC;
mem[16'h0D52] = 8'hDC;
mem[16'h0D53] = 8'hDC;
mem[16'h0D54] = 8'hDC;
mem[16'h0D55] = 8'hDC;
mem[16'h0D56] = 8'hDC;
mem[16'h0D57] = 8'hDC;
mem[16'h0D58] = 8'hDC;
mem[16'h0D59] = 8'hDC;
mem[16'h0D5A] = 8'hDC;
mem[16'h0D5B] = 8'hDC;
mem[16'h0D5C] = 8'hDC;
mem[16'h0D5D] = 8'hDC;
mem[16'h0D5E] = 8'hDC;
mem[16'h0D5F] = 8'hDC;
mem[16'h0D60] = 8'hDC;
mem[16'h0D61] = 8'hDC;
mem[16'h0D62] = 8'hDC;
mem[16'h0D63] = 8'hDC;
mem[16'h0D64] = 8'hDC;
mem[16'h0D65] = 8'hDC;
mem[16'h0D66] = 8'hDC;
mem[16'h0D67] = 8'hDC;
mem[16'h0D68] = 8'hDC;
mem[16'h0D69] = 8'hDC;
mem[16'h0D6A] = 8'hDC;
mem[16'h0D6B] = 8'hDC;
mem[16'h0D6C] = 8'hDC;
mem[16'h0D6D] = 8'hDC;
mem[16'h0D6E] = 8'hDC;
mem[16'h0D6F] = 8'hDC;
mem[16'h0D70] = 8'hDC;
mem[16'h0D71] = 8'hDC;
mem[16'h0D72] = 8'hDC;
mem[16'h0D73] = 8'hDC;
mem[16'h0D74] = 8'hDC;
mem[16'h0D75] = 8'hDC;
mem[16'h0D76] = 8'hDC;
mem[16'h0D77] = 8'hDC;
mem[16'h0D78] = 8'hDC;
mem[16'h0D79] = 8'hDC;
mem[16'h0D7A] = 8'hDC;
mem[16'h0D7B] = 8'hDC;
mem[16'h0D7C] = 8'hDC;
mem[16'h0D7D] = 8'hDC;
mem[16'h0D7E] = 8'hDC;
mem[16'h0D7F] = 8'hDC;
mem[16'h0D80] = 8'hDC;
mem[16'h0D81] = 8'hDC;
mem[16'h0D82] = 8'hDC;
mem[16'h0D83] = 8'hDC;
mem[16'h0D84] = 8'hDC;
mem[16'h0D85] = 8'hDC;
mem[16'h0D86] = 8'hDC;
mem[16'h0D87] = 8'hDC;
mem[16'h0D88] = 8'hDC;
mem[16'h0D89] = 8'hDC;
mem[16'h0D8A] = 8'hDC;
mem[16'h0D8B] = 8'hDC;
mem[16'h0D8C] = 8'hDC;
mem[16'h0D8D] = 8'hDC;
mem[16'h0D8E] = 8'hDC;
mem[16'h0D8F] = 8'hDC;
mem[16'h0D90] = 8'hDC;
mem[16'h0D91] = 8'hDC;
mem[16'h0D92] = 8'hDC;
mem[16'h0D93] = 8'hDC;
mem[16'h0D94] = 8'hDC;
mem[16'h0D95] = 8'hDC;
mem[16'h0D96] = 8'hDC;
mem[16'h0D97] = 8'hDC;
mem[16'h0D98] = 8'hDC;
mem[16'h0D99] = 8'hDC;
mem[16'h0D9A] = 8'hDC;
mem[16'h0D9B] = 8'hDC;
mem[16'h0D9C] = 8'hDC;
mem[16'h0D9D] = 8'hDC;
mem[16'h0D9E] = 8'hDC;
mem[16'h0D9F] = 8'hDC;
mem[16'h0DA0] = 8'hDC;
mem[16'h0DA1] = 8'hDC;
mem[16'h0DA2] = 8'hDC;
mem[16'h0DA3] = 8'hDC;
mem[16'h0DA4] = 8'hDC;
mem[16'h0DA5] = 8'hDC;
mem[16'h0DA6] = 8'hDC;
mem[16'h0DA7] = 8'hDC;
mem[16'h0DA8] = 8'hDC;
mem[16'h0DA9] = 8'hDC;
mem[16'h0DAA] = 8'hDC;
mem[16'h0DAB] = 8'hDC;
mem[16'h0DAC] = 8'hDC;
mem[16'h0DAD] = 8'hDC;
mem[16'h0DAE] = 8'hDC;
mem[16'h0DAF] = 8'hDC;
mem[16'h0DB0] = 8'hDC;
mem[16'h0DB1] = 8'hDC;
mem[16'h0DB2] = 8'hDC;
mem[16'h0DB3] = 8'hDC;
mem[16'h0DB4] = 8'hDC;
mem[16'h0DB5] = 8'hDC;
mem[16'h0DB6] = 8'hDC;
mem[16'h0DB7] = 8'hDC;
mem[16'h0DB8] = 8'hDC;
mem[16'h0DB9] = 8'hDC;
mem[16'h0DBA] = 8'hDC;
mem[16'h0DBB] = 8'hDC;
mem[16'h0DBC] = 8'hDC;
mem[16'h0DBD] = 8'hDC;
mem[16'h0DBE] = 8'hDC;
mem[16'h0DBF] = 8'hDC;
mem[16'h0DC0] = 8'hDC;
mem[16'h0DC1] = 8'hDC;
mem[16'h0DC2] = 8'hDC;
mem[16'h0DC3] = 8'hDC;
mem[16'h0DC4] = 8'hDC;
mem[16'h0DC5] = 8'hDC;
mem[16'h0DC6] = 8'hDC;
mem[16'h0DC7] = 8'hDC;
mem[16'h0DC8] = 8'hDC;
mem[16'h0DC9] = 8'hDC;
mem[16'h0DCA] = 8'hDC;
mem[16'h0DCB] = 8'hDC;
mem[16'h0DCC] = 8'hDC;
mem[16'h0DCD] = 8'hDC;
mem[16'h0DCE] = 8'hDC;
mem[16'h0DCF] = 8'hDC;
mem[16'h0DD0] = 8'hDC;
mem[16'h0DD1] = 8'hDC;
mem[16'h0DD2] = 8'hDC;
mem[16'h0DD3] = 8'hDC;
mem[16'h0DD4] = 8'hDC;
mem[16'h0DD5] = 8'hDC;
mem[16'h0DD6] = 8'hDC;
mem[16'h0DD7] = 8'hDC;
mem[16'h0DD8] = 8'hDC;
mem[16'h0DD9] = 8'hDC;
mem[16'h0DDA] = 8'hDC;
mem[16'h0DDB] = 8'hDC;
mem[16'h0DDC] = 8'hDC;
mem[16'h0DDD] = 8'hDC;
mem[16'h0DDE] = 8'hDC;
mem[16'h0DDF] = 8'hDC;
mem[16'h0DE0] = 8'hDC;
mem[16'h0DE1] = 8'hDC;
mem[16'h0DE2] = 8'hDC;
mem[16'h0DE3] = 8'hDC;
mem[16'h0DE4] = 8'hDC;
mem[16'h0DE5] = 8'hDC;
mem[16'h0DE6] = 8'hDC;
mem[16'h0DE7] = 8'hDC;
mem[16'h0DE8] = 8'hDC;
mem[16'h0DE9] = 8'hDC;
mem[16'h0DEA] = 8'hDC;
mem[16'h0DEB] = 8'hDC;
mem[16'h0DEC] = 8'hDC;
mem[16'h0DED] = 8'hDC;
mem[16'h0DEE] = 8'hDC;
mem[16'h0DEF] = 8'hDC;
mem[16'h0DF0] = 8'hDC;
mem[16'h0DF1] = 8'hDC;
mem[16'h0DF2] = 8'hDC;
mem[16'h0DF3] = 8'hDC;
mem[16'h0DF4] = 8'hDC;
mem[16'h0DF5] = 8'hDC;
mem[16'h0DF6] = 8'hDC;
mem[16'h0DF7] = 8'hDC;
mem[16'h0DF8] = 8'hDC;
mem[16'h0DF9] = 8'hDC;
mem[16'h0DFA] = 8'hDC;
mem[16'h0DFB] = 8'hDC;
mem[16'h0DFC] = 8'hDC;
mem[16'h0DFD] = 8'hDC;
mem[16'h0DFE] = 8'hDC;
mem[16'h0DFF] = 8'hDC;
mem[16'h0E00] = 8'h00;
mem[16'h0E01] = 8'h9C;
mem[16'h0E02] = 8'h00;
mem[16'h0E03] = 8'h08;
mem[16'h0E04] = 8'h3A;
mem[16'h0E05] = 8'h03;
mem[16'h0E06] = 8'h00;
mem[16'h0E07] = 8'h00;
mem[16'h0E08] = 8'h00;
mem[16'h0E09] = 8'hC0;
mem[16'h0E0A] = 8'h60;
mem[16'h0E0B] = 8'h01;
mem[16'h0E0C] = 8'h05;
mem[16'h0E0D] = 8'h00;
mem[16'h0E0E] = 8'h00;
mem[16'h0E0F] = 8'h6B;
mem[16'h0E10] = 8'h00;
mem[16'h0E11] = 8'h9C;
mem[16'h0E12] = 8'h00;
mem[16'h0E13] = 8'h04;
mem[16'h0E14] = 8'h00;
mem[16'h0E15] = 8'h00;
mem[16'h0E16] = 8'h00;
mem[16'h0E17] = 8'h00;
mem[16'h0E18] = 8'hFF;
mem[16'h0E19] = 8'h0C;
mem[16'h0E1A] = 8'h00;
mem[16'h0E1B] = 8'h56;
mem[16'h0E1C] = 8'hFF;
mem[16'h0E1D] = 8'hFF;
mem[16'h0E1E] = 8'h00;
mem[16'h0E1F] = 8'h00;
mem[16'h0E20] = 8'h00;
mem[16'h0E21] = 8'h28;
mem[16'h0E22] = 8'h00;
mem[16'h0E23] = 8'h18;
mem[16'h0E24] = 8'h00;
mem[16'h0E25] = 8'h01;
mem[16'h0E26] = 8'h00;
mem[16'h0E27] = 8'h09;
mem[16'h0E28] = 8'h80;
mem[16'h0E29] = 8'h04;
mem[16'h0E2A] = 8'hD0;
mem[16'h0E2B] = 8'h07;
mem[16'h0E2C] = 8'h00;
mem[16'h0E2D] = 8'h00;
mem[16'h0E2E] = 8'hE8;
mem[16'h0E2F] = 8'h01;
mem[16'h0E30] = 8'hFE;
mem[16'h0E31] = 8'h00;
mem[16'h0E32] = 8'hFF;
mem[16'h0E33] = 8'hAA;
mem[16'h0E34] = 8'h05;
mem[16'h0E35] = 8'h28;
mem[16'h0E36] = 8'h09;
mem[16'h0E37] = 8'h03;
mem[16'h0E38] = 8'h1B;
mem[16'h0E39] = 8'hFD;
mem[16'h0E3A] = 8'h00;
mem[16'h0E3B] = 8'h9C;
mem[16'h0E3C] = 8'h00;
mem[16'h0E3D] = 8'h9C;
mem[16'h0E3E] = 8'h00;
mem[16'h0E3F] = 8'h9C;
mem[16'h0E40] = 8'h00;
mem[16'h0E41] = 8'h9C;
mem[16'h0E42] = 8'hA2;
mem[16'h0E43] = 8'h5B;
mem[16'h0E44] = 8'h82;
mem[16'h0E45] = 8'h98;
mem[16'h0E46] = 8'h62;
mem[16'h0E47] = 8'hD8;
mem[16'h0E48] = 8'h00;
mem[16'h0E49] = 8'hB7;
mem[16'h0E4A] = 8'h00;
mem[16'h0E4B] = 8'h00;
mem[16'h0E4C] = 8'hFF;
mem[16'h0E4D] = 8'hFF;
mem[16'h0E4E] = 8'h4E;
mem[16'h0E4F] = 8'h6E;
mem[16'h0E50] = 8'h69;
mem[16'h0E51] = 8'hFF;
mem[16'h0E52] = 8'h55;
mem[16'h0E53] = 8'h52;
mem[16'h0E54] = 8'h00;
mem[16'h0E55] = 8'h28;
mem[16'h0E56] = 8'h61;
mem[16'h0E57] = 8'h08;
mem[16'h0E58] = 8'hFF;
mem[16'h0E59] = 8'hFF;
mem[16'h0E5A] = 8'h00;
mem[16'h0E5B] = 8'h00;
mem[16'h0E5C] = 8'hFF;
mem[16'h0E5D] = 8'hFF;
mem[16'h0E5E] = 8'h38;
mem[16'h0E5F] = 8'hDE;
mem[16'h0E60] = 8'hA5;
mem[16'h0E61] = 8'h00;
mem[16'h0E62] = 8'h00;
mem[16'h0E63] = 8'h00;
mem[16'h0E64] = 8'hFF;
mem[16'h0E65] = 8'hFF;
mem[16'h0E66] = 8'h00;
mem[16'h0E67] = 8'h01;
mem[16'h0E68] = 8'h08;
mem[16'h0E69] = 8'h04;
mem[16'h0E6A] = 8'h08;
mem[16'h0E6B] = 8'h04;
mem[16'h0E6C] = 8'h08;
mem[16'h0E6D] = 8'h04;
mem[16'h0E6E] = 8'h08;
mem[16'h0E6F] = 8'h00;
mem[16'h0E70] = 8'h96;
mem[16'h0E71] = 8'hFF;
mem[16'h0E72] = 8'h00;
mem[16'h0E73] = 8'h00;
mem[16'h0E74] = 8'h96;
mem[16'h0E75] = 8'h18;
mem[16'h0E76] = 8'hFF;
mem[16'h0E77] = 8'h18;
mem[16'h0E78] = 8'h01;
mem[16'h0E79] = 8'h16;
mem[16'h0E7A] = 8'h00;
mem[16'h0E7B] = 8'h00;
mem[16'h0E7C] = 8'hFF;
mem[16'h0E7D] = 8'hC1;
mem[16'h0E7E] = 8'hDA;
mem[16'h0E7F] = 8'h88;
mem[16'h0E80] = 8'h95;
mem[16'h0E81] = 8'hFF;
mem[16'h0E82] = 8'h00;
mem[16'h0E83] = 8'h00;
mem[16'h0E84] = 8'hFF;
mem[16'h0E85] = 8'h00;
mem[16'h0E86] = 8'h00;
mem[16'h0E87] = 8'hFF;
mem[16'h0E88] = 8'hFF;
mem[16'h0E89] = 8'h00;
mem[16'h0E8A] = 8'h00;
mem[16'h0E8B] = 8'h00;
mem[16'h0E8C] = 8'hFF;
mem[16'h0E8D] = 8'hFF;
mem[16'h0E8E] = 8'h00;
mem[16'h0E8F] = 8'h03;
mem[16'h0E90] = 8'h4C;
mem[16'h0E91] = 8'h64;
mem[16'h0E92] = 8'h00;
mem[16'h0E93] = 8'h00;
mem[16'h0E94] = 8'hFF;
mem[16'h0E95] = 8'hFF;
mem[16'h0E96] = 8'h00;
mem[16'h0E97] = 8'h00;
mem[16'h0E98] = 8'hFF;
mem[16'h0E99] = 8'h00;
mem[16'h0E9A] = 8'h00;
mem[16'h0E9B] = 8'h00;
mem[16'h0E9C] = 8'h00;
mem[16'h0E9D] = 8'h88;
mem[16'h0E9E] = 8'hFF;
mem[16'h0E9F] = 8'hFF;
mem[16'h0EA0] = 8'hFF;
mem[16'h0EA1] = 8'h69;
mem[16'h0EA2] = 8'hFF;
mem[16'h0EA3] = 8'h00;
mem[16'h0EA4] = 8'h00;
mem[16'h0EA5] = 8'hD0;
mem[16'h0EA6] = 8'hD1;
mem[16'h0EA7] = 8'hFF;
mem[16'h0EA8] = 8'hFF;
mem[16'h0EA9] = 8'h69;
mem[16'h0EAA] = 8'hFF;
mem[16'h0EAB] = 8'hFF;
mem[16'h0EAC] = 8'h00;
mem[16'h0EAD] = 8'h09;
mem[16'h0EAE] = 8'h08;
mem[16'h0EAF] = 8'h04;
mem[16'h0EB0] = 8'h08;
mem[16'h0EB1] = 8'hE6;
mem[16'h0EB2] = 8'hB8;
mem[16'h0EB3] = 8'hD0;
mem[16'h0EB4] = 8'h02;
mem[16'h0EB5] = 8'hE6;
mem[16'h0EB6] = 8'hB9;
mem[16'h0EB7] = 8'hAD;
mem[16'h0EB8] = 8'h05;
mem[16'h0EB9] = 8'h02;
mem[16'h0EBA] = 8'hC9;
mem[16'h0EBB] = 8'h3A;
mem[16'h0EBC] = 8'hB0;
mem[16'h0EBD] = 8'h0A;
mem[16'h0EBE] = 8'hC9;
mem[16'h0EBF] = 8'h20;
mem[16'h0EC0] = 8'hF0;
mem[16'h0EC1] = 8'hEF;
mem[16'h0EC2] = 8'h38;
mem[16'h0EC3] = 8'hE9;
mem[16'h0EC4] = 8'h30;
mem[16'h0EC5] = 8'h38;
mem[16'h0EC6] = 8'hE9;
mem[16'h0EC7] = 8'hD0;
mem[16'h0EC8] = 8'h60;
mem[16'h0EC9] = 8'h80;
mem[16'h0ECA] = 8'h4F;
mem[16'h0ECB] = 8'hC7;
mem[16'h0ECC] = 8'h52;
mem[16'h0ECD] = 8'hFF;
mem[16'h0ECE] = 8'h00;
mem[16'h0ECF] = 8'h00;
mem[16'h0ED0] = 8'hFF;
mem[16'h0ED1] = 8'hFF;
mem[16'h0ED2] = 8'h00;
mem[16'h0ED3] = 8'h00;
mem[16'h0ED4] = 8'hFF;
mem[16'h0ED5] = 8'hFF;
mem[16'h0ED6] = 8'h00;
mem[16'h0ED7] = 8'h00;
mem[16'h0ED8] = 8'h00;
mem[16'h0ED9] = 8'hFF;
mem[16'h0EDA] = 8'h00;
mem[16'h0EDB] = 8'h00;
mem[16'h0EDC] = 8'hFF;
mem[16'h0EDD] = 8'hFF;
mem[16'h0EDE] = 8'h00;
mem[16'h0EDF] = 8'h00;
mem[16'h0EE0] = 8'hFF;
mem[16'h0EE1] = 8'hFF;
mem[16'h0EE2] = 8'h00;
mem[16'h0EE3] = 8'h00;
mem[16'h0EE4] = 8'hFF;
mem[16'h0EE5] = 8'hFF;
mem[16'h0EE6] = 8'h00;
mem[16'h0EE7] = 8'h00;
mem[16'h0EE8] = 8'hFF;
mem[16'h0EE9] = 8'hFF;
mem[16'h0EEA] = 8'h00;
mem[16'h0EEB] = 8'h00;
mem[16'h0EEC] = 8'hFF;
mem[16'h0EED] = 8'hFF;
mem[16'h0EEE] = 8'h00;
mem[16'h0EEF] = 8'h00;
mem[16'h0EF0] = 8'hFF;
mem[16'h0EF1] = 8'h01;
mem[16'h0EF2] = 8'h00;
mem[16'h0EF3] = 8'h00;
mem[16'h0EF4] = 8'hFF;
mem[16'h0EF5] = 8'hFF;
mem[16'h0EF6] = 8'h00;
mem[16'h0EF7] = 8'h00;
mem[16'h0EF8] = 8'hF8;
mem[16'h0EF9] = 8'hFF;
mem[16'h0EFA] = 8'h00;
mem[16'h0EFB] = 8'h00;
mem[16'h0EFC] = 8'hFF;
mem[16'h0EFD] = 8'hFF;
mem[16'h0EFE] = 8'h00;
mem[16'h0EFF] = 8'h10;
mem[16'h0F00] = 8'h00;
mem[16'h0F01] = 8'hFF;
mem[16'h0F02] = 8'h00;
mem[16'h0F03] = 8'h00;
mem[16'h0F04] = 8'h00;
mem[16'h0F05] = 8'hFF;
mem[16'h0F06] = 8'h00;
mem[16'h0F07] = 8'h00;
mem[16'h0F08] = 8'h00;
mem[16'h0F09] = 8'hFF;
mem[16'h0F0A] = 8'h00;
mem[16'h0F0B] = 8'h00;
mem[16'h0F0C] = 8'h00;
mem[16'h0F0D] = 8'hFF;
mem[16'h0F0E] = 8'h00;
mem[16'h0F0F] = 8'h00;
mem[16'h0F10] = 8'h00;
mem[16'h0F11] = 8'hFF;
mem[16'h0F12] = 8'h00;
mem[16'h0F13] = 8'h00;
mem[16'h0F14] = 8'h00;
mem[16'h0F15] = 8'hFF;
mem[16'h0F16] = 8'h00;
mem[16'h0F17] = 8'h00;
mem[16'h0F18] = 8'h00;
mem[16'h0F19] = 8'hFF;
mem[16'h0F1A] = 8'h00;
mem[16'h0F1B] = 8'h00;
mem[16'h0F1C] = 8'h00;
mem[16'h0F1D] = 8'hFF;
mem[16'h0F1E] = 8'h00;
mem[16'h0F1F] = 8'h00;
mem[16'h0F20] = 8'h00;
mem[16'h0F21] = 8'hFF;
mem[16'h0F22] = 8'h00;
mem[16'h0F23] = 8'h00;
mem[16'h0F24] = 8'h00;
mem[16'h0F25] = 8'hFF;
mem[16'h0F26] = 8'h00;
mem[16'h0F27] = 8'h00;
mem[16'h0F28] = 8'h00;
mem[16'h0F29] = 8'hFF;
mem[16'h0F2A] = 8'h00;
mem[16'h0F2B] = 8'h00;
mem[16'h0F2C] = 8'h00;
mem[16'h0F2D] = 8'hFF;
mem[16'h0F2E] = 8'h00;
mem[16'h0F2F] = 8'h00;
mem[16'h0F30] = 8'h00;
mem[16'h0F31] = 8'hFF;
mem[16'h0F32] = 8'h00;
mem[16'h0F33] = 8'h00;
mem[16'h0F34] = 8'h00;
mem[16'h0F35] = 8'hFF;
mem[16'h0F36] = 8'h00;
mem[16'h0F37] = 8'h00;
mem[16'h0F38] = 8'h00;
mem[16'h0F39] = 8'hFF;
mem[16'h0F3A] = 8'h00;
mem[16'h0F3B] = 8'h00;
mem[16'h0F3C] = 8'h00;
mem[16'h0F3D] = 8'hFF;
mem[16'h0F3E] = 8'h00;
mem[16'h0F3F] = 8'h00;
mem[16'h0F40] = 8'h00;
mem[16'h0F41] = 8'hFF;
mem[16'h0F42] = 8'h00;
mem[16'h0F43] = 8'h00;
mem[16'h0F44] = 8'h00;
mem[16'h0F45] = 8'hFF;
mem[16'h0F46] = 8'h00;
mem[16'h0F47] = 8'h00;
mem[16'h0F48] = 8'h00;
mem[16'h0F49] = 8'hFF;
mem[16'h0F4A] = 8'h00;
mem[16'h0F4B] = 8'h00;
mem[16'h0F4C] = 8'h00;
mem[16'h0F4D] = 8'hFF;
mem[16'h0F4E] = 8'h00;
mem[16'h0F4F] = 8'h00;
mem[16'h0F50] = 8'h00;
mem[16'h0F51] = 8'hFF;
mem[16'h0F52] = 8'h00;
mem[16'h0F53] = 8'h00;
mem[16'h0F54] = 8'h00;
mem[16'h0F55] = 8'hFF;
mem[16'h0F56] = 8'h00;
mem[16'h0F57] = 8'h00;
mem[16'h0F58] = 8'h00;
mem[16'h0F59] = 8'hFF;
mem[16'h0F5A] = 8'h00;
mem[16'h0F5B] = 8'h00;
mem[16'h0F5C] = 8'h00;
mem[16'h0F5D] = 8'hFF;
mem[16'h0F5E] = 8'h00;
mem[16'h0F5F] = 8'h00;
mem[16'h0F60] = 8'h00;
mem[16'h0F61] = 8'hFF;
mem[16'h0F62] = 8'h00;
mem[16'h0F63] = 8'h00;
mem[16'h0F64] = 8'h00;
mem[16'h0F65] = 8'hFF;
mem[16'h0F66] = 8'h00;
mem[16'h0F67] = 8'h00;
mem[16'h0F68] = 8'h00;
mem[16'h0F69] = 8'hFF;
mem[16'h0F6A] = 8'h00;
mem[16'h0F6B] = 8'h00;
mem[16'h0F6C] = 8'h00;
mem[16'h0F6D] = 8'hFF;
mem[16'h0F6E] = 8'h00;
mem[16'h0F6F] = 8'h00;
mem[16'h0F70] = 8'h00;
mem[16'h0F71] = 8'hFF;
mem[16'h0F72] = 8'h00;
mem[16'h0F73] = 8'h00;
mem[16'h0F74] = 8'h00;
mem[16'h0F75] = 8'hFF;
mem[16'h0F76] = 8'h00;
mem[16'h0F77] = 8'h00;
mem[16'h0F78] = 8'h00;
mem[16'h0F79] = 8'hFF;
mem[16'h0F7A] = 8'h00;
mem[16'h0F7B] = 8'h00;
mem[16'h0F7C] = 8'h00;
mem[16'h0F7D] = 8'hFF;
mem[16'h0F7E] = 8'h00;
mem[16'h0F7F] = 8'h00;
mem[16'h0F80] = 8'h00;
mem[16'h0F81] = 8'hFF;
mem[16'h0F82] = 8'h00;
mem[16'h0F83] = 8'h00;
mem[16'h0F84] = 8'h00;
mem[16'h0F85] = 8'hFF;
mem[16'h0F86] = 8'h00;
mem[16'h0F87] = 8'h00;
mem[16'h0F88] = 8'h00;
mem[16'h0F89] = 8'hFF;
mem[16'h0F8A] = 8'h00;
mem[16'h0F8B] = 8'h00;
mem[16'h0F8C] = 8'h00;
mem[16'h0F8D] = 8'hFF;
mem[16'h0F8E] = 8'h00;
mem[16'h0F8F] = 8'h00;
mem[16'h0F90] = 8'h00;
mem[16'h0F91] = 8'hFF;
mem[16'h0F92] = 8'h00;
mem[16'h0F93] = 8'h00;
mem[16'h0F94] = 8'h00;
mem[16'h0F95] = 8'hFF;
mem[16'h0F96] = 8'h00;
mem[16'h0F97] = 8'h00;
mem[16'h0F98] = 8'h00;
mem[16'h0F99] = 8'hFF;
mem[16'h0F9A] = 8'h00;
mem[16'h0F9B] = 8'h00;
mem[16'h0F9C] = 8'h00;
mem[16'h0F9D] = 8'hFF;
mem[16'h0F9E] = 8'h00;
mem[16'h0F9F] = 8'h00;
mem[16'h0FA0] = 8'h00;
mem[16'h0FA1] = 8'hFF;
mem[16'h0FA2] = 8'h00;
mem[16'h0FA3] = 8'h00;
mem[16'h0FA4] = 8'h00;
mem[16'h0FA5] = 8'hFF;
mem[16'h0FA6] = 8'h00;
mem[16'h0FA7] = 8'h00;
mem[16'h0FA8] = 8'h00;
mem[16'h0FA9] = 8'hFF;
mem[16'h0FAA] = 8'h00;
mem[16'h0FAB] = 8'h00;
mem[16'h0FAC] = 8'h00;
mem[16'h0FAD] = 8'hFF;
mem[16'h0FAE] = 8'h00;
mem[16'h0FAF] = 8'h00;
mem[16'h0FB0] = 8'h00;
mem[16'h0FB1] = 8'hFF;
mem[16'h0FB2] = 8'h00;
mem[16'h0FB3] = 8'h00;
mem[16'h0FB4] = 8'h00;
mem[16'h0FB5] = 8'hFF;
mem[16'h0FB6] = 8'h00;
mem[16'h0FB7] = 8'h00;
mem[16'h0FB8] = 8'h00;
mem[16'h0FB9] = 8'hFF;
mem[16'h0FBA] = 8'h00;
mem[16'h0FBB] = 8'h00;
mem[16'h0FBC] = 8'h00;
mem[16'h0FBD] = 8'hFF;
mem[16'h0FBE] = 8'h00;
mem[16'h0FBF] = 8'h00;
mem[16'h0FC0] = 8'h00;
mem[16'h0FC1] = 8'hFF;
mem[16'h0FC2] = 8'h00;
mem[16'h0FC3] = 8'h00;
mem[16'h0FC4] = 8'h00;
mem[16'h0FC5] = 8'hFF;
mem[16'h0FC6] = 8'h00;
mem[16'h0FC7] = 8'h00;
mem[16'h0FC8] = 8'h00;
mem[16'h0FC9] = 8'hFF;
mem[16'h0FCA] = 8'h39;
mem[16'h0FCB] = 8'hB5;
mem[16'h0FCC] = 8'h38;
mem[16'h0FCD] = 8'hB7;
mem[16'h0FCE] = 8'hDA;
mem[16'h0FCF] = 8'hB6;
mem[16'h0FD0] = 8'h4F;
mem[16'h0FD1] = 8'hB6;
mem[16'h0FD2] = 8'h5F;
mem[16'h0FD3] = 8'hBF;
mem[16'h0FD4] = 8'h20;
mem[16'h0FD5] = 8'hB4;
mem[16'h0FD6] = 8'h09;
mem[16'h0FD7] = 8'h00;
mem[16'h0FD8] = 8'hB0;
mem[16'h0FD9] = 8'h02;
mem[16'h0FDA] = 8'h10;
mem[16'h0FDB] = 8'hCF;
mem[16'h0FDC] = 8'h5F;
mem[16'h0FDD] = 8'h0B;
mem[16'h0FDE] = 8'h40;
mem[16'h0FDF] = 8'h84;
mem[16'h0FE0] = 8'hFF;
mem[16'h0FE1] = 8'h26;
mem[16'h0FE2] = 8'hFC;
mem[16'h0FE3] = 8'hA0;
mem[16'h0FE4] = 8'h37;
mem[16'h0FE5] = 8'hFD;
mem[16'h0FE6] = 8'h77;
mem[16'h0FE7] = 8'hFD;
mem[16'h0FE8] = 8'h9B;
mem[16'h0FE9] = 8'hF5;
mem[16'h0FEA] = 8'h84;
mem[16'h0FEB] = 8'hFF;
mem[16'h0FEC] = 8'hB5;
mem[16'h0FED] = 8'h3B;
mem[16'h0FEE] = 8'h9C;
mem[16'h0FEF] = 8'hCF;
mem[16'h0FF0] = 8'h5F;
mem[16'h0FF1] = 8'h0B;
mem[16'h0FF2] = 8'h40;
mem[16'h0FF3] = 8'h69;
mem[16'h0FF4] = 8'h00;
mem[16'h0FF5] = 8'h6F;
mem[16'h0FF6] = 8'h00;
mem[16'h0FF7] = 8'h22;
mem[16'h0FF8] = 8'h00;
mem[16'h0FF9] = 8'hC1;
mem[16'h0FFA] = 8'h00;
mem[16'h0FFB] = 8'h00;
mem[16'h0FFC] = 8'h00;
mem[16'h0FFD] = 8'h01;
mem[16'h0FFE] = 8'h00;
mem[16'h0FFF] = 8'h37;
mem[16'h1000] = 8'hB9;
mem[16'h1001] = 8'hC3;
mem[16'h1002] = 8'hB0;
mem[16'h1003] = 8'hB0;
mem[16'h1004] = 8'hC7;
mem[16'h1005] = 8'h8D;
mem[16'h1006] = 8'hC6;
mem[16'h1007] = 8'hB5;
mem[16'h1008] = 8'hB9;
mem[16'h1009] = 8'h8D;
mem[16'h100A] = 8'hD8;
mem[16'h100B] = 8'h8D;
mem[16'h100C] = 8'h8D;
mem[16'h100D] = 8'hB1;
mem[16'h100E] = 8'h8D;
mem[16'h100F] = 8'hAC;
mem[16'h1010] = 8'h00;
mem[16'h1011] = 8'hA4;
mem[16'h1012] = 8'h00;
mem[16'h1013] = 8'hB0;
mem[16'h1014] = 8'h00;
mem[16'h1015] = 8'hB0;
mem[16'h1016] = 8'h00;
mem[16'h1017] = 8'hCC;
mem[16'h1018] = 8'h00;
mem[16'h1019] = 8'hB2;
mem[16'h101A] = 8'h00;
mem[16'h101B] = 8'hB0;
mem[16'h101C] = 8'h00;
mem[16'h101D] = 8'h8D;
mem[16'h101E] = 8'h00;
mem[16'h101F] = 8'h00;
mem[16'h1020] = 8'h00;
mem[16'h1021] = 8'hFF;
mem[16'h1022] = 8'h00;
mem[16'h1023] = 8'h02;
mem[16'h1024] = 8'h00;
mem[16'h1025] = 8'hFF;
mem[16'h1026] = 8'h00;
mem[16'h1027] = 8'h02;
mem[16'h1028] = 8'h00;
mem[16'h1029] = 8'hFF;
mem[16'h102A] = 8'h00;
mem[16'h102B] = 8'h02;
mem[16'h102C] = 8'h00;
mem[16'h102D] = 8'hFF;
mem[16'h102E] = 8'h00;
mem[16'h102F] = 8'h02;
mem[16'h1030] = 8'h00;
mem[16'h1031] = 8'hFF;
mem[16'h1032] = 8'h00;
mem[16'h1033] = 8'h00;
mem[16'h1034] = 8'h00;
mem[16'h1035] = 8'hFF;
mem[16'h1036] = 8'h00;
mem[16'h1037] = 8'h00;
mem[16'h1038] = 8'h00;
mem[16'h1039] = 8'hFF;
mem[16'h103A] = 8'h00;
mem[16'h103B] = 8'h00;
mem[16'h103C] = 8'h00;
mem[16'h103D] = 8'hFF;
mem[16'h103E] = 8'h00;
mem[16'h103F] = 8'h00;
mem[16'h1040] = 8'h00;
mem[16'h1041] = 8'hFF;
mem[16'h1042] = 8'h00;
mem[16'h1043] = 8'h00;
mem[16'h1044] = 8'h00;
mem[16'h1045] = 8'hFF;
mem[16'h1046] = 8'h00;
mem[16'h1047] = 8'h00;
mem[16'h1048] = 8'h00;
mem[16'h1049] = 8'hFF;
mem[16'h104A] = 8'h00;
mem[16'h104B] = 8'h00;
mem[16'h104C] = 8'h00;
mem[16'h104D] = 8'hFF;
mem[16'h104E] = 8'h00;
mem[16'h104F] = 8'h00;
mem[16'h1050] = 8'h00;
mem[16'h1051] = 8'hFF;
mem[16'h1052] = 8'h00;
mem[16'h1053] = 8'h00;
mem[16'h1054] = 8'h00;
mem[16'h1055] = 8'hFF;
mem[16'h1056] = 8'h00;
mem[16'h1057] = 8'h00;
mem[16'h1058] = 8'h00;
mem[16'h1059] = 8'hFF;
mem[16'h105A] = 8'h00;
mem[16'h105B] = 8'h00;
mem[16'h105C] = 8'h00;
mem[16'h105D] = 8'hFF;
mem[16'h105E] = 8'h00;
mem[16'h105F] = 8'h00;
mem[16'h1060] = 8'h00;
mem[16'h1061] = 8'hFF;
mem[16'h1062] = 8'h00;
mem[16'h1063] = 8'h00;
mem[16'h1064] = 8'h00;
mem[16'h1065] = 8'hFF;
mem[16'h1066] = 8'h00;
mem[16'h1067] = 8'h00;
mem[16'h1068] = 8'h00;
mem[16'h1069] = 8'hFF;
mem[16'h106A] = 8'h00;
mem[16'h106B] = 8'h00;
mem[16'h106C] = 8'h00;
mem[16'h106D] = 8'hFF;
mem[16'h106E] = 8'h00;
mem[16'h106F] = 8'h00;
mem[16'h1070] = 8'h00;
mem[16'h1071] = 8'hFF;
mem[16'h1072] = 8'h00;
mem[16'h1073] = 8'h00;
mem[16'h1074] = 8'h00;
mem[16'h1075] = 8'hFF;
mem[16'h1076] = 8'h00;
mem[16'h1077] = 8'h00;
mem[16'h1078] = 8'h00;
mem[16'h1079] = 8'hFF;
mem[16'h107A] = 8'h00;
mem[16'h107B] = 8'h00;
mem[16'h107C] = 8'h00;
mem[16'h107D] = 8'hFF;
mem[16'h107E] = 8'h00;
mem[16'h107F] = 8'h00;
mem[16'h1080] = 8'h00;
mem[16'h1081] = 8'hFF;
mem[16'h1082] = 8'h00;
mem[16'h1083] = 8'h00;
mem[16'h1084] = 8'h00;
mem[16'h1085] = 8'hFF;
mem[16'h1086] = 8'h00;
mem[16'h1087] = 8'h00;
mem[16'h1088] = 8'h00;
mem[16'h1089] = 8'hFF;
mem[16'h108A] = 8'h00;
mem[16'h108B] = 8'h00;
mem[16'h108C] = 8'h00;
mem[16'h108D] = 8'hFF;
mem[16'h108E] = 8'h00;
mem[16'h108F] = 8'h02;
mem[16'h1090] = 8'h00;
mem[16'h1091] = 8'hFF;
mem[16'h1092] = 8'h00;
mem[16'h1093] = 8'h00;
mem[16'h1094] = 8'h00;
mem[16'h1095] = 8'hFF;
mem[16'h1096] = 8'h00;
mem[16'h1097] = 8'h00;
mem[16'h1098] = 8'h00;
mem[16'h1099] = 8'hFF;
mem[16'h109A] = 8'h00;
mem[16'h109B] = 8'h00;
mem[16'h109C] = 8'h00;
mem[16'h109D] = 8'hFF;
mem[16'h109E] = 8'h00;
mem[16'h109F] = 8'h00;
mem[16'h10A0] = 8'h00;
mem[16'h10A1] = 8'hFF;
mem[16'h10A2] = 8'h00;
mem[16'h10A3] = 8'h02;
mem[16'h10A4] = 8'h00;
mem[16'h10A5] = 8'hFF;
mem[16'h10A6] = 8'h00;
mem[16'h10A7] = 8'h02;
mem[16'h10A8] = 8'h00;
mem[16'h10A9] = 8'hFF;
mem[16'h10AA] = 8'h00;
mem[16'h10AB] = 8'h00;
mem[16'h10AC] = 8'h00;
mem[16'h10AD] = 8'hFF;
mem[16'h10AE] = 8'h00;
mem[16'h10AF] = 8'h02;
mem[16'h10B0] = 8'h00;
mem[16'h10B1] = 8'hFF;
mem[16'h10B2] = 8'h00;
mem[16'h10B3] = 8'h00;
mem[16'h10B4] = 8'h00;
mem[16'h10B5] = 8'hFF;
mem[16'h10B6] = 8'h00;
mem[16'h10B7] = 8'h00;
mem[16'h10B8] = 8'h00;
mem[16'h10B9] = 8'hFF;
mem[16'h10BA] = 8'h00;
mem[16'h10BB] = 8'h00;
mem[16'h10BC] = 8'h00;
mem[16'h10BD] = 8'hFF;
mem[16'h10BE] = 8'h00;
mem[16'h10BF] = 8'h00;
mem[16'h10C0] = 8'h00;
mem[16'h10C1] = 8'hFF;
mem[16'h10C2] = 8'h00;
mem[16'h10C3] = 8'h00;
mem[16'h10C4] = 8'h00;
mem[16'h10C5] = 8'hFF;
mem[16'h10C6] = 8'h00;
mem[16'h10C7] = 8'h00;
mem[16'h10C8] = 8'h00;
mem[16'h10C9] = 8'hFF;
mem[16'h10CA] = 8'h00;
mem[16'h10CB] = 8'h00;
mem[16'h10CC] = 8'h00;
mem[16'h10CD] = 8'hFF;
mem[16'h10CE] = 8'h00;
mem[16'h10CF] = 8'h00;
mem[16'h10D0] = 8'h00;
mem[16'h10D1] = 8'hFF;
mem[16'h10D2] = 8'h00;
mem[16'h10D3] = 8'h00;
mem[16'h10D4] = 8'h00;
mem[16'h10D5] = 8'hFF;
mem[16'h10D6] = 8'h00;
mem[16'h10D7] = 8'h00;
mem[16'h10D8] = 8'h00;
mem[16'h10D9] = 8'hFF;
mem[16'h10DA] = 8'h00;
mem[16'h10DB] = 8'h00;
mem[16'h10DC] = 8'h00;
mem[16'h10DD] = 8'hFF;
mem[16'h10DE] = 8'h00;
mem[16'h10DF] = 8'h00;
mem[16'h10E0] = 8'h00;
mem[16'h10E1] = 8'hFF;
mem[16'h10E2] = 8'h00;
mem[16'h10E3] = 8'h00;
mem[16'h10E4] = 8'h00;
mem[16'h10E5] = 8'hFF;
mem[16'h10E6] = 8'h00;
mem[16'h10E7] = 8'h00;
mem[16'h10E8] = 8'h00;
mem[16'h10E9] = 8'hFF;
mem[16'h10EA] = 8'h00;
mem[16'h10EB] = 8'h00;
mem[16'h10EC] = 8'h00;
mem[16'h10ED] = 8'hFF;
mem[16'h10EE] = 8'h00;
mem[16'h10EF] = 8'h00;
mem[16'h10F0] = 8'h00;
mem[16'h10F1] = 8'hFF;
mem[16'h10F2] = 8'h00;
mem[16'h10F3] = 8'h00;
mem[16'h10F4] = 8'h00;
mem[16'h10F5] = 8'hFF;
mem[16'h10F6] = 8'h00;
mem[16'h10F7] = 8'h00;
mem[16'h10F8] = 8'h00;
mem[16'h10F9] = 8'hFF;
mem[16'h10FA] = 8'h00;
mem[16'h10FB] = 8'h00;
mem[16'h10FC] = 8'h00;
mem[16'h10FD] = 8'hFF;
mem[16'h10FE] = 8'h00;
mem[16'h10FF] = 8'h00;
mem[16'h1100] = 8'hA0;
mem[16'h1101] = 8'h03;
mem[16'h1102] = 8'h84;
mem[16'h1103] = 8'h37;
mem[16'h1104] = 8'hA0;
mem[16'h1105] = 8'h09;
mem[16'h1106] = 8'h84;
mem[16'h1107] = 8'h36;
mem[16'h1108] = 8'h60;
mem[16'h1109] = 8'h48;
mem[16'h110A] = 8'h84;
mem[16'h110B] = 8'h4E;
mem[16'h110C] = 8'hC9;
mem[16'h110D] = 8'h8D;
mem[16'h110E] = 8'hF0;
mem[16'h110F] = 8'h68;
mem[16'h1110] = 8'hA5;
mem[16'h1111] = 8'h25;
mem[16'h1112] = 8'h4A;
mem[16'h1113] = 8'h29;
mem[16'h1114] = 8'h03;
mem[16'h1115] = 8'h09;
mem[16'h1116] = 8'h20;
mem[16'h1117] = 8'h85;
mem[16'h1118] = 8'h2B;
mem[16'h1119] = 8'hA5;
mem[16'h111A] = 8'h25;
mem[16'h111B] = 8'h6A;
mem[16'h111C] = 8'h08;
mem[16'h111D] = 8'h0A;
mem[16'h111E] = 8'h29;
mem[16'h111F] = 8'h18;
mem[16'h1120] = 8'h85;
mem[16'h1121] = 8'h2A;
mem[16'h1122] = 8'h0A;
mem[16'h1123] = 8'h0A;
mem[16'h1124] = 8'h05;
mem[16'h1125] = 8'h2A;
mem[16'h1126] = 8'h0A;
mem[16'h1127] = 8'h28;
mem[16'h1128] = 8'h6A;
mem[16'h1129] = 8'h18;
mem[16'h112A] = 8'h65;
mem[16'h112B] = 8'h24;
mem[16'h112C] = 8'h85;
mem[16'h112D] = 8'h2A;
mem[16'h112E] = 8'h68;
mem[16'h112F] = 8'h29;
mem[16'h1130] = 8'h7F;
mem[16'h1131] = 8'h48;
mem[16'h1132] = 8'hA9;
mem[16'h1133] = 8'h00;
mem[16'h1134] = 8'h85;
mem[16'h1135] = 8'h27;
mem[16'h1136] = 8'h68;
mem[16'h1137] = 8'h48;
mem[16'h1138] = 8'h2A;
mem[16'h1139] = 8'h26;
mem[16'h113A] = 8'h27;
mem[16'h113B] = 8'h2A;
mem[16'h113C] = 8'h26;
mem[16'h113D] = 8'h27;
mem[16'h113E] = 8'h2A;
mem[16'h113F] = 8'h26;
mem[16'h1140] = 8'h27;
mem[16'h1141] = 8'h85;
mem[16'h1142] = 8'h26;
mem[16'h1143] = 8'hA5;
mem[16'h1144] = 8'h27;
mem[16'h1145] = 8'h18;
mem[16'h1146] = 8'h69;
mem[16'h1147] = 8'h04;
mem[16'h1148] = 8'h85;
mem[16'h1149] = 8'h27;
mem[16'h114A] = 8'hA0;
mem[16'h114B] = 8'h00;
mem[16'h114C] = 8'hB1;
mem[16'h114D] = 8'h26;
mem[16'h114E] = 8'h48;
mem[16'h114F] = 8'h84;
mem[16'h1150] = 8'h4F;
mem[16'h1151] = 8'hA0;
mem[16'h1152] = 8'h00;
mem[16'h1153] = 8'h51;
mem[16'h1154] = 8'h2A;
mem[16'h1155] = 8'h91;
mem[16'h1156] = 8'h2A;
mem[16'h1157] = 8'hA5;
mem[16'h1158] = 8'h2B;
mem[16'h1159] = 8'hEA;
mem[16'h115A] = 8'hEA;
mem[16'h115B] = 8'h85;
mem[16'h115C] = 8'h2B;
mem[16'h115D] = 8'h68;
mem[16'h115E] = 8'h51;
mem[16'h115F] = 8'h2A;
mem[16'h1160] = 8'hEA;
mem[16'h1161] = 8'hEA;
mem[16'h1162] = 8'hA4;
mem[16'h1163] = 8'h4F;
mem[16'h1164] = 8'hA5;
mem[16'h1165] = 8'h2B;
mem[16'h1166] = 8'h18;
mem[16'h1167] = 8'h69;
mem[16'h1168] = 8'h04;
mem[16'h1169] = 8'h85;
mem[16'h116A] = 8'h2B;
mem[16'h116B] = 8'hC8;
mem[16'h116C] = 8'hC0;
mem[16'h116D] = 8'h08;
mem[16'h116E] = 8'hD0;
mem[16'h116F] = 8'hDC;
mem[16'h1170] = 8'hE6;
mem[16'h1171] = 8'h24;
mem[16'h1172] = 8'hA5;
mem[16'h1173] = 8'h24;
mem[16'h1174] = 8'hC5;
mem[16'h1175] = 8'h21;
mem[16'h1176] = 8'h90;
mem[16'h1177] = 8'h10;
mem[16'h1178] = 8'hA5;
mem[16'h1179] = 8'h20;
mem[16'h117A] = 8'h85;
mem[16'h117B] = 8'h24;
mem[16'h117C] = 8'hE6;
mem[16'h117D] = 8'h25;
mem[16'h117E] = 8'hA5;
mem[16'h117F] = 8'h25;
mem[16'h1180] = 8'hC5;
mem[16'h1181] = 8'h23;
mem[16'h1182] = 8'h90;
mem[16'h1183] = 8'h04;
mem[16'h1184] = 8'hA5;
mem[16'h1185] = 8'h22;
mem[16'h1186] = 8'h85;
mem[16'h1187] = 8'h25;
mem[16'h1188] = 8'hA4;
mem[16'h1189] = 8'h4E;
mem[16'h118A] = 8'h68;
mem[16'h118B] = 8'h60;
mem[16'h118C] = 8'hFF;
mem[16'h118D] = 8'hFF;
mem[16'h118E] = 8'h00;
mem[16'h118F] = 8'h00;
mem[16'h1190] = 8'hFF;
mem[16'h1191] = 8'hFF;
mem[16'h1192] = 8'h00;
mem[16'h1193] = 8'h00;
mem[16'h1194] = 8'hFF;
mem[16'h1195] = 8'hFF;
mem[16'h1196] = 8'h00;
mem[16'h1197] = 8'h00;
mem[16'h1198] = 8'hFF;
mem[16'h1199] = 8'hFF;
mem[16'h119A] = 8'h00;
mem[16'h119B] = 8'h00;
mem[16'h119C] = 8'hFF;
mem[16'h119D] = 8'hFF;
mem[16'h119E] = 8'h00;
mem[16'h119F] = 8'h00;
mem[16'h11A0] = 8'hFF;
mem[16'h11A1] = 8'hFF;
mem[16'h11A2] = 8'h00;
mem[16'h11A3] = 8'h00;
mem[16'h11A4] = 8'hFF;
mem[16'h11A5] = 8'hFF;
mem[16'h11A6] = 8'h00;
mem[16'h11A7] = 8'h00;
mem[16'h11A8] = 8'hFF;
mem[16'h11A9] = 8'hFF;
mem[16'h11AA] = 8'h00;
mem[16'h11AB] = 8'h00;
mem[16'h11AC] = 8'hFF;
mem[16'h11AD] = 8'hFF;
mem[16'h11AE] = 8'h00;
mem[16'h11AF] = 8'h00;
mem[16'h11B0] = 8'hFF;
mem[16'h11B1] = 8'hFF;
mem[16'h11B2] = 8'h00;
mem[16'h11B3] = 8'h00;
mem[16'h11B4] = 8'hFF;
mem[16'h11B5] = 8'hFF;
mem[16'h11B6] = 8'h00;
mem[16'h11B7] = 8'h00;
mem[16'h11B8] = 8'hFF;
mem[16'h11B9] = 8'hFF;
mem[16'h11BA] = 8'h00;
mem[16'h11BB] = 8'h00;
mem[16'h11BC] = 8'hFF;
mem[16'h11BD] = 8'hFF;
mem[16'h11BE] = 8'h00;
mem[16'h11BF] = 8'h00;
mem[16'h11C0] = 8'h00;
mem[16'h11C1] = 8'h00;
mem[16'h11C2] = 8'h00;
mem[16'h11C3] = 8'h00;
mem[16'h11C4] = 8'h00;
mem[16'h11C5] = 8'h00;
mem[16'h11C6] = 8'h00;
mem[16'h11C7] = 8'h00;
mem[16'h11C8] = 8'h00;
mem[16'h11C9] = 8'h00;
mem[16'h11CA] = 8'h00;
mem[16'h11CB] = 8'h00;
mem[16'h11CC] = 8'hB6;
mem[16'h11CD] = 8'h00;
mem[16'h11CE] = 8'h00;
mem[16'h11CF] = 8'h00;
mem[16'h11D0] = 8'h4C;
mem[16'h11D1] = 8'hBF;
mem[16'h11D2] = 8'h9D;
mem[16'h11D3] = 8'h4C;
mem[16'h11D4] = 8'h84;
mem[16'h11D5] = 8'h9D;
mem[16'h11D6] = 8'h4C;
mem[16'h11D7] = 8'hFD;
mem[16'h11D8] = 8'hAA;
mem[16'h11D9] = 8'h4C;
mem[16'h11DA] = 8'hB5;
mem[16'h11DB] = 8'hB7;
mem[16'h11DC] = 8'hAD;
mem[16'h11DD] = 8'h0F;
mem[16'h11DE] = 8'h9D;
mem[16'h11DF] = 8'hAC;
mem[16'h11E0] = 8'h0E;
mem[16'h11E1] = 8'h9D;
mem[16'h11E2] = 8'h60;
mem[16'h11E3] = 8'hAD;
mem[16'h11E4] = 8'hC2;
mem[16'h11E5] = 8'hAA;
mem[16'h11E6] = 8'hAC;
mem[16'h11E7] = 8'hC1;
mem[16'h11E8] = 8'hAA;
mem[16'h11E9] = 8'h60;
mem[16'h11EA] = 8'h4C;
mem[16'h11EB] = 8'h51;
mem[16'h11EC] = 8'hA8;
mem[16'h11ED] = 8'hEA;
mem[16'h11EE] = 8'hEA;
mem[16'h11EF] = 8'h4C;
mem[16'h11F0] = 8'h59;
mem[16'h11F1] = 8'hFA;
mem[16'h11F2] = 8'h43;
mem[16'h11F3] = 8'h00;
mem[16'h11F4] = 8'h95;
mem[16'h11F5] = 8'h4C;
mem[16'h11F6] = 8'h58;
mem[16'h11F7] = 8'hFF;
mem[16'h11F8] = 8'h4C;
mem[16'h11F9] = 8'h65;
mem[16'h11FA] = 8'hFF;
mem[16'h11FB] = 8'h4C;
mem[16'h11FC] = 8'h65;
mem[16'h11FD] = 8'hFF;
mem[16'h11FE] = 8'h65;
mem[16'h11FF] = 8'hFF;
mem[16'h1200] = 8'h00;
mem[16'h1201] = 8'hFF;
mem[16'h1202] = 8'hFF;
mem[16'h1203] = 8'h00;
mem[16'h1204] = 8'h00;
mem[16'h1205] = 8'hFF;
mem[16'h1206] = 8'hFF;
mem[16'h1207] = 8'h00;
mem[16'h1208] = 8'h00;
mem[16'h1209] = 8'hFF;
mem[16'h120A] = 8'hFF;
mem[16'h120B] = 8'h00;
mem[16'h120C] = 8'h00;
mem[16'h120D] = 8'hFF;
mem[16'h120E] = 8'hFF;
mem[16'h120F] = 8'h00;
mem[16'h1210] = 8'h00;
mem[16'h1211] = 8'hFF;
mem[16'h1212] = 8'hFF;
mem[16'h1213] = 8'h00;
mem[16'h1214] = 8'h00;
mem[16'h1215] = 8'hFF;
mem[16'h1216] = 8'hFF;
mem[16'h1217] = 8'h00;
mem[16'h1218] = 8'h00;
mem[16'h1219] = 8'hFF;
mem[16'h121A] = 8'hFF;
mem[16'h121B] = 8'h00;
mem[16'h121C] = 8'h00;
mem[16'h121D] = 8'hFF;
mem[16'h121E] = 8'hFF;
mem[16'h121F] = 8'h00;
mem[16'h1220] = 8'h00;
mem[16'h1221] = 8'hFF;
mem[16'h1222] = 8'hFF;
mem[16'h1223] = 8'h00;
mem[16'h1224] = 8'h00;
mem[16'h1225] = 8'hFF;
mem[16'h1226] = 8'hFF;
mem[16'h1227] = 8'h00;
mem[16'h1228] = 8'h00;
mem[16'h1229] = 8'hFF;
mem[16'h122A] = 8'hFF;
mem[16'h122B] = 8'h00;
mem[16'h122C] = 8'h00;
mem[16'h122D] = 8'hFF;
mem[16'h122E] = 8'hFF;
mem[16'h122F] = 8'h00;
mem[16'h1230] = 8'h00;
mem[16'h1231] = 8'hFF;
mem[16'h1232] = 8'hFF;
mem[16'h1233] = 8'h00;
mem[16'h1234] = 8'h00;
mem[16'h1235] = 8'hFF;
mem[16'h1236] = 8'hFF;
mem[16'h1237] = 8'h00;
mem[16'h1238] = 8'h00;
mem[16'h1239] = 8'h14;
mem[16'h123A] = 8'h22;
mem[16'h123B] = 8'h22;
mem[16'h123C] = 8'h22;
mem[16'h123D] = 8'h41;
mem[16'h123E] = 8'h7F;
mem[16'h123F] = 8'h08;
mem[16'h1240] = 8'h10;
mem[16'h1241] = 8'h08;
mem[16'h1242] = 8'h04;
mem[16'h1243] = 8'h7E;
mem[16'h1244] = 8'h04;
mem[16'h1245] = 8'h08;
mem[16'h1246] = 8'h10;
mem[16'h1247] = 8'h00;
mem[16'h1248] = 8'h08;
mem[16'h1249] = 8'h10;
mem[16'h124A] = 8'h20;
mem[16'h124B] = 8'h7E;
mem[16'h124C] = 8'h20;
mem[16'h124D] = 8'h10;
mem[16'h124E] = 8'h08;
mem[16'h124F] = 8'h00;
mem[16'h1250] = 8'h08;
mem[16'h1251] = 8'h08;
mem[16'h1252] = 8'h08;
mem[16'h1253] = 8'h49;
mem[16'h1254] = 8'h2A;
mem[16'h1255] = 8'h1C;
mem[16'h1256] = 8'h08;
mem[16'h1257] = 8'h00;
mem[16'h1258] = 8'h08;
mem[16'h1259] = 8'h1C;
mem[16'h125A] = 8'h2A;
mem[16'h125B] = 8'h49;
mem[16'h125C] = 8'h08;
mem[16'h125D] = 8'h08;
mem[16'h125E] = 8'h08;
mem[16'h125F] = 8'h00;
mem[16'h1260] = 8'h08;
mem[16'h1261] = 8'h49;
mem[16'h1262] = 8'h2A;
mem[16'h1263] = 8'h1C;
mem[16'h1264] = 8'h49;
mem[16'h1265] = 8'h2A;
mem[16'h1266] = 8'h1C;
mem[16'h1267] = 8'h08;
mem[16'h1268] = 8'h40;
mem[16'h1269] = 8'h60;
mem[16'h126A] = 8'h70;
mem[16'h126B] = 8'h78;
mem[16'h126C] = 8'h70;
mem[16'h126D] = 8'h60;
mem[16'h126E] = 8'h40;
mem[16'h126F] = 8'h00;
mem[16'h1270] = 8'h40;
mem[16'h1271] = 8'h40;
mem[16'h1272] = 8'h20;
mem[16'h1273] = 8'h20;
mem[16'h1274] = 8'h13;
mem[16'h1275] = 8'h14;
mem[16'h1276] = 8'h0C;
mem[16'h1277] = 8'h08;
mem[16'h1278] = 8'h1A;
mem[16'h1279] = 8'h00;
mem[16'h127A] = 8'h00;
mem[16'h127B] = 8'h7C;
mem[16'h127C] = 8'h2A;
mem[16'h127D] = 8'h28;
mem[16'h127E] = 8'h34;
mem[16'h127F] = 8'h00;
mem[16'h1280] = 8'h36;
mem[16'h1281] = 8'h7F;
mem[16'h1282] = 8'h7F;
mem[16'h1283] = 8'h7F;
mem[16'h1284] = 8'h3E;
mem[16'h1285] = 8'h1C;
mem[16'h1286] = 8'h08;
mem[16'h1287] = 8'h00;
mem[16'h1288] = 8'h08;
mem[16'h1289] = 8'h1C;
mem[16'h128A] = 8'h3E;
mem[16'h128B] = 8'h7F;
mem[16'h128C] = 8'h3E;
mem[16'h128D] = 8'h1C;
mem[16'h128E] = 8'h08;
mem[16'h128F] = 8'h00;
mem[16'h1290] = 8'h08;
mem[16'h1291] = 8'h1C;
mem[16'h1292] = 8'h3E;
mem[16'h1293] = 8'h7F;
mem[16'h1294] = 8'h7F;
mem[16'h1295] = 8'h2A;
mem[16'h1296] = 8'h08;
mem[16'h1297] = 8'h00;
mem[16'h1298] = 8'h08;
mem[16'h1299] = 8'h1C;
mem[16'h129A] = 8'h1C;
mem[16'h129B] = 8'h2A;
mem[16'h129C] = 8'h7F;
mem[16'h129D] = 8'h7F;
mem[16'h129E] = 8'h2A;
mem[16'h129F] = 8'h08;
mem[16'h12A0] = 8'h3E;
mem[16'h12A1] = 8'h08;
mem[16'h12A2] = 8'h08;
mem[16'h12A3] = 8'h22;
mem[16'h12A4] = 8'h36;
mem[16'h12A5] = 8'h2A;
mem[16'h12A6] = 8'h22;
mem[16'h12A7] = 8'h00;
mem[16'h12A8] = 8'h00;
mem[16'h12A9] = 8'h22;
mem[16'h12AA] = 8'h14;
mem[16'h12AB] = 8'h08;
mem[16'h12AC] = 8'h14;
mem[16'h12AD] = 8'h22;
mem[16'h12AE] = 8'h00;
mem[16'h12AF] = 8'h00;
mem[16'h12B0] = 8'h04;
mem[16'h12B1] = 8'h0E;
mem[16'h12B2] = 8'h04;
mem[16'h12B3] = 8'h04;
mem[16'h12B4] = 8'h00;
mem[16'h12B5] = 8'h00;
mem[16'h12B6] = 8'h00;
mem[16'h12B7] = 8'h00;
mem[16'h12B8] = 8'h00;
mem[16'h12B9] = 8'h08;
mem[16'h12BA] = 8'h00;
mem[16'h12BB] = 8'h3E;
mem[16'h12BC] = 8'h00;
mem[16'h12BD] = 8'h08;
mem[16'h12BE] = 8'h00;
mem[16'h12BF] = 8'h00;
mem[16'h12C0] = 8'h18;
mem[16'h12C1] = 8'h24;
mem[16'h12C2] = 8'h08;
mem[16'h12C3] = 8'h14;
mem[16'h12C4] = 8'h08;
mem[16'h12C5] = 8'h12;
mem[16'h12C6] = 8'h0C;
mem[16'h12C7] = 8'h00;
mem[16'h12C8] = 8'h10;
mem[16'h12C9] = 8'h38;
mem[16'h12CA] = 8'h04;
mem[16'h12CB] = 8'h04;
mem[16'h12CC] = 8'h38;
mem[16'h12CD] = 8'h10;
mem[16'h12CE] = 8'h00;
mem[16'h12CF] = 8'h00;
mem[16'h12D0] = 8'h08;
mem[16'h12D1] = 8'h1C;
mem[16'h12D2] = 8'h08;
mem[16'h12D3] = 8'h1C;
mem[16'h12D4] = 8'h3E;
mem[16'h12D5] = 8'h1C;
mem[16'h12D6] = 8'h3E;
mem[16'h12D7] = 8'h7F;
mem[16'h12D8] = 8'h08;
mem[16'h12D9] = 8'h3E;
mem[16'h12DA] = 8'h1C;
mem[16'h12DB] = 8'h08;
mem[16'h12DC] = 8'h1C;
mem[16'h12DD] = 8'h1C;
mem[16'h12DE] = 8'h3E;
mem[16'h12DF] = 8'h7F;
mem[16'h12E0] = 8'h00;
mem[16'h12E1] = 8'h2A;
mem[16'h12E2] = 8'h3E;
mem[16'h12E3] = 8'h1C;
mem[16'h12E4] = 8'h1C;
mem[16'h12E5] = 8'h1C;
mem[16'h12E6] = 8'h3E;
mem[16'h12E7] = 8'h7F;
mem[16'h12E8] = 8'h00;
mem[16'h12E9] = 8'h10;
mem[16'h12EA] = 8'h3C;
mem[16'h12EB] = 8'h3E;
mem[16'h12EC] = 8'h18;
mem[16'h12ED] = 8'h0C;
mem[16'h12EE] = 8'h1E;
mem[16'h12EF] = 8'h3F;
mem[16'h12F0] = 8'h00;
mem[16'h12F1] = 8'h08;
mem[16'h12F2] = 8'h18;
mem[16'h12F3] = 8'h3A;
mem[16'h12F4] = 8'h7B;
mem[16'h12F5] = 8'h3E;
mem[16'h12F6] = 8'h1C;
mem[16'h12F7] = 8'h7F;
mem[16'h12F8] = 8'h04;
mem[16'h12F9] = 8'h00;
mem[16'h12FA] = 8'h08;
mem[16'h12FB] = 8'h1C;
mem[16'h12FC] = 8'h1C;
mem[16'h12FD] = 8'h08;
mem[16'h12FE] = 8'h1C;
mem[16'h12FF] = 8'h3E;
mem[16'h1300] = 8'h00;
mem[16'h1301] = 8'h00;
mem[16'h1302] = 8'h00;
mem[16'h1303] = 8'h00;
mem[16'h1304] = 8'h00;
mem[16'h1305] = 8'h00;
mem[16'h1306] = 8'h00;
mem[16'h1307] = 8'h00;
mem[16'h1308] = 8'h10;
mem[16'h1309] = 8'h10;
mem[16'h130A] = 8'h10;
mem[16'h130B] = 8'h10;
mem[16'h130C] = 8'h00;
mem[16'h130D] = 8'h00;
mem[16'h130E] = 8'h10;
mem[16'h130F] = 8'h00;
mem[16'h1310] = 8'h24;
mem[16'h1311] = 8'h24;
mem[16'h1312] = 8'h24;
mem[16'h1313] = 8'h00;
mem[16'h1314] = 8'h00;
mem[16'h1315] = 8'h00;
mem[16'h1316] = 8'h00;
mem[16'h1317] = 8'h00;
mem[16'h1318] = 8'h24;
mem[16'h1319] = 8'h24;
mem[16'h131A] = 8'h7E;
mem[16'h131B] = 8'h24;
mem[16'h131C] = 8'h7E;
mem[16'h131D] = 8'h24;
mem[16'h131E] = 8'h24;
mem[16'h131F] = 8'h00;
mem[16'h1320] = 8'h10;
mem[16'h1321] = 8'h78;
mem[16'h1322] = 8'h14;
mem[16'h1323] = 8'h38;
mem[16'h1324] = 8'h50;
mem[16'h1325] = 8'h3C;
mem[16'h1326] = 8'h10;
mem[16'h1327] = 8'h00;
mem[16'h1328] = 8'h00;
mem[16'h1329] = 8'h46;
mem[16'h132A] = 8'h26;
mem[16'h132B] = 8'h10;
mem[16'h132C] = 8'h08;
mem[16'h132D] = 8'h64;
mem[16'h132E] = 8'h62;
mem[16'h132F] = 8'h00;
mem[16'h1330] = 8'h0C;
mem[16'h1331] = 8'h12;
mem[16'h1332] = 8'h12;
mem[16'h1333] = 8'h0C;
mem[16'h1334] = 8'h52;
mem[16'h1335] = 8'h22;
mem[16'h1336] = 8'h5C;
mem[16'h1337] = 8'h00;
mem[16'h1338] = 8'h20;
mem[16'h1339] = 8'h10;
mem[16'h133A] = 8'h08;
mem[16'h133B] = 8'h00;
mem[16'h133C] = 8'h00;
mem[16'h133D] = 8'h00;
mem[16'h133E] = 8'h00;
mem[16'h133F] = 8'h00;
mem[16'h1340] = 8'h20;
mem[16'h1341] = 8'h10;
mem[16'h1342] = 8'h08;
mem[16'h1343] = 8'h08;
mem[16'h1344] = 8'h08;
mem[16'h1345] = 8'h10;
mem[16'h1346] = 8'h20;
mem[16'h1347] = 8'h00;
mem[16'h1348] = 8'h04;
mem[16'h1349] = 8'h08;
mem[16'h134A] = 8'h10;
mem[16'h134B] = 8'h10;
mem[16'h134C] = 8'h10;
mem[16'h134D] = 8'h08;
mem[16'h134E] = 8'h04;
mem[16'h134F] = 8'h00;
mem[16'h1350] = 8'h10;
mem[16'h1351] = 8'h54;
mem[16'h1352] = 8'h38;
mem[16'h1353] = 8'h7C;
mem[16'h1354] = 8'h38;
mem[16'h1355] = 8'h54;
mem[16'h1356] = 8'h10;
mem[16'h1357] = 8'h00;
mem[16'h1358] = 8'h00;
mem[16'h1359] = 8'h10;
mem[16'h135A] = 8'h10;
mem[16'h135B] = 8'h7C;
mem[16'h135C] = 8'h10;
mem[16'h135D] = 8'h10;
mem[16'h135E] = 8'h00;
mem[16'h135F] = 8'h00;
mem[16'h1360] = 8'h00;
mem[16'h1361] = 8'h00;
mem[16'h1362] = 8'h00;
mem[16'h1363] = 8'h00;
mem[16'h1364] = 8'h00;
mem[16'h1365] = 8'h18;
mem[16'h1366] = 8'h18;
mem[16'h1367] = 8'h0C;
mem[16'h1368] = 8'h00;
mem[16'h1369] = 8'h00;
mem[16'h136A] = 8'h00;
mem[16'h136B] = 8'h7E;
mem[16'h136C] = 8'h00;
mem[16'h136D] = 8'h00;
mem[16'h136E] = 8'h00;
mem[16'h136F] = 8'h00;
mem[16'h1370] = 8'h00;
mem[16'h1371] = 8'h00;
mem[16'h1372] = 8'h00;
mem[16'h1373] = 8'h00;
mem[16'h1374] = 8'h00;
mem[16'h1375] = 8'h18;
mem[16'h1376] = 8'h18;
mem[16'h1377] = 8'h00;
mem[16'h1378] = 8'h28;
mem[16'h1379] = 8'h40;
mem[16'h137A] = 8'h20;
mem[16'h137B] = 8'h10;
mem[16'h137C] = 8'h08;
mem[16'h137D] = 8'h04;
mem[16'h137E] = 8'h02;
mem[16'h137F] = 8'h00;
mem[16'h1380] = 8'h3C;
mem[16'h1381] = 8'h42;
mem[16'h1382] = 8'h42;
mem[16'h1383] = 8'h42;
mem[16'h1384] = 8'h42;
mem[16'h1385] = 8'h42;
mem[16'h1386] = 8'h3C;
mem[16'h1387] = 8'h00;
mem[16'h1388] = 8'h10;
mem[16'h1389] = 8'h18;
mem[16'h138A] = 8'h14;
mem[16'h138B] = 8'h10;
mem[16'h138C] = 8'h10;
mem[16'h138D] = 8'h10;
mem[16'h138E] = 8'h7C;
mem[16'h138F] = 8'h00;
mem[16'h1390] = 8'h3C;
mem[16'h1391] = 8'h42;
mem[16'h1392] = 8'h40;
mem[16'h1393] = 8'h30;
mem[16'h1394] = 8'h0C;
mem[16'h1395] = 8'h02;
mem[16'h1396] = 8'h7E;
mem[16'h1397] = 8'h00;
mem[16'h1398] = 8'h3C;
mem[16'h1399] = 8'h42;
mem[16'h139A] = 8'h40;
mem[16'h139B] = 8'h38;
mem[16'h139C] = 8'h40;
mem[16'h139D] = 8'h42;
mem[16'h139E] = 8'h3C;
mem[16'h139F] = 8'h00;
mem[16'h13A0] = 8'h20;
mem[16'h13A1] = 8'h30;
mem[16'h13A2] = 8'h28;
mem[16'h13A3] = 8'h24;
mem[16'h13A4] = 8'h7E;
mem[16'h13A5] = 8'h20;
mem[16'h13A6] = 8'h20;
mem[16'h13A7] = 8'h00;
mem[16'h13A8] = 8'h7E;
mem[16'h13A9] = 8'h02;
mem[16'h13AA] = 8'h1E;
mem[16'h13AB] = 8'h20;
mem[16'h13AC] = 8'h40;
mem[16'h13AD] = 8'h22;
mem[16'h13AE] = 8'h1C;
mem[16'h13AF] = 8'h00;
mem[16'h13B0] = 8'h38;
mem[16'h13B1] = 8'h04;
mem[16'h13B2] = 8'h02;
mem[16'h13B3] = 8'h3E;
mem[16'h13B4] = 8'h42;
mem[16'h13B5] = 8'h42;
mem[16'h13B6] = 8'h3C;
mem[16'h13B7] = 8'h00;
mem[16'h13B8] = 8'h7E;
mem[16'h13B9] = 8'h42;
mem[16'h13BA] = 8'h20;
mem[16'h13BB] = 8'h10;
mem[16'h13BC] = 8'h08;
mem[16'h13BD] = 8'h08;
mem[16'h13BE] = 8'h08;
mem[16'h13BF] = 8'h00;
mem[16'h13C0] = 8'h3C;
mem[16'h13C1] = 8'h42;
mem[16'h13C2] = 8'h42;
mem[16'h13C3] = 8'h3C;
mem[16'h13C4] = 8'h42;
mem[16'h13C5] = 8'h42;
mem[16'h13C6] = 8'h3C;
mem[16'h13C7] = 8'h00;
mem[16'h13C8] = 8'h3C;
mem[16'h13C9] = 8'h42;
mem[16'h13CA] = 8'h42;
mem[16'h13CB] = 8'h7C;
mem[16'h13CC] = 8'h40;
mem[16'h13CD] = 8'h20;
mem[16'h13CE] = 8'h1C;
mem[16'h13CF] = 8'h00;
mem[16'h13D0] = 8'h00;
mem[16'h13D1] = 8'h00;
mem[16'h13D2] = 8'h18;
mem[16'h13D3] = 8'h18;
mem[16'h13D4] = 8'h00;
mem[16'h13D5] = 8'h18;
mem[16'h13D6] = 8'h18;
mem[16'h13D7] = 8'h00;
mem[16'h13D8] = 8'h00;
mem[16'h13D9] = 8'h00;
mem[16'h13DA] = 8'h18;
mem[16'h13DB] = 8'h18;
mem[16'h13DC] = 8'h00;
mem[16'h13DD] = 8'h18;
mem[16'h13DE] = 8'h18;
mem[16'h13DF] = 8'h0C;
mem[16'h13E0] = 8'h20;
mem[16'h13E1] = 8'h10;
mem[16'h13E2] = 8'h08;
mem[16'h13E3] = 8'h04;
mem[16'h13E4] = 8'h08;
mem[16'h13E5] = 8'h10;
mem[16'h13E6] = 8'h20;
mem[16'h13E7] = 8'h00;
mem[16'h13E8] = 8'h00;
mem[16'h13E9] = 8'h00;
mem[16'h13EA] = 8'h3E;
mem[16'h13EB] = 8'h00;
mem[16'h13EC] = 8'h3E;
mem[16'h13ED] = 8'h00;
mem[16'h13EE] = 8'h00;
mem[16'h13EF] = 8'h00;
mem[16'h13F0] = 8'h04;
mem[16'h13F1] = 8'h08;
mem[16'h13F2] = 8'h10;
mem[16'h13F3] = 8'h20;
mem[16'h13F4] = 8'h10;
mem[16'h13F5] = 8'h08;
mem[16'h13F6] = 8'h04;
mem[16'h13F7] = 8'h00;
mem[16'h13F8] = 8'h60;
mem[16'h13F9] = 8'h42;
mem[16'h13FA] = 8'h40;
mem[16'h13FB] = 8'h30;
mem[16'h13FC] = 8'h08;
mem[16'h13FD] = 8'h00;
mem[16'h13FE] = 8'h08;
mem[16'h13FF] = 8'h00;
mem[16'h1400] = 8'h38;
mem[16'h1401] = 8'h44;
mem[16'h1402] = 8'h52;
mem[16'h1403] = 8'h6A;
mem[16'h1404] = 8'h32;
mem[16'h1405] = 8'h04;
mem[16'h1406] = 8'h78;
mem[16'h1407] = 8'h00;
mem[16'h1408] = 8'h18;
mem[16'h1409] = 8'h24;
mem[16'h140A] = 8'h42;
mem[16'h140B] = 8'h7E;
mem[16'h140C] = 8'h42;
mem[16'h140D] = 8'h42;
mem[16'h140E] = 8'h42;
mem[16'h140F] = 8'h00;
mem[16'h1410] = 8'h3E;
mem[16'h1411] = 8'h44;
mem[16'h1412] = 8'h44;
mem[16'h1413] = 8'h3C;
mem[16'h1414] = 8'h44;
mem[16'h1415] = 8'h44;
mem[16'h1416] = 8'h3E;
mem[16'h1417] = 8'h00;
mem[16'h1418] = 8'h3C;
mem[16'h1419] = 8'h42;
mem[16'h141A] = 8'h02;
mem[16'h141B] = 8'h02;
mem[16'h141C] = 8'h02;
mem[16'h141D] = 8'h42;
mem[16'h141E] = 8'h3C;
mem[16'h141F] = 8'h00;
mem[16'h1420] = 8'h3E;
mem[16'h1421] = 8'h44;
mem[16'h1422] = 8'h44;
mem[16'h1423] = 8'h44;
mem[16'h1424] = 8'h44;
mem[16'h1425] = 8'h44;
mem[16'h1426] = 8'h3E;
mem[16'h1427] = 8'h00;
mem[16'h1428] = 8'h7E;
mem[16'h1429] = 8'h02;
mem[16'h142A] = 8'h02;
mem[16'h142B] = 8'h1E;
mem[16'h142C] = 8'h02;
mem[16'h142D] = 8'h02;
mem[16'h142E] = 8'h7E;
mem[16'h142F] = 8'h00;
mem[16'h1430] = 8'h7E;
mem[16'h1431] = 8'h02;
mem[16'h1432] = 8'h02;
mem[16'h1433] = 8'h1E;
mem[16'h1434] = 8'h02;
mem[16'h1435] = 8'h02;
mem[16'h1436] = 8'h02;
mem[16'h1437] = 8'h00;
mem[16'h1438] = 8'h3C;
mem[16'h1439] = 8'h42;
mem[16'h143A] = 8'h02;
mem[16'h143B] = 8'h72;
mem[16'h143C] = 8'h42;
mem[16'h143D] = 8'h42;
mem[16'h143E] = 8'h3C;
mem[16'h143F] = 8'h00;
mem[16'h1440] = 8'h42;
mem[16'h1441] = 8'h42;
mem[16'h1442] = 8'h42;
mem[16'h1443] = 8'h7E;
mem[16'h1444] = 8'h42;
mem[16'h1445] = 8'h42;
mem[16'h1446] = 8'h42;
mem[16'h1447] = 8'h00;
mem[16'h1448] = 8'h38;
mem[16'h1449] = 8'h10;
mem[16'h144A] = 8'h10;
mem[16'h144B] = 8'h10;
mem[16'h144C] = 8'h10;
mem[16'h144D] = 8'h10;
mem[16'h144E] = 8'h38;
mem[16'h144F] = 8'h00;
mem[16'h1450] = 8'h70;
mem[16'h1451] = 8'h20;
mem[16'h1452] = 8'h20;
mem[16'h1453] = 8'h20;
mem[16'h1454] = 8'h20;
mem[16'h1455] = 8'h22;
mem[16'h1456] = 8'h1C;
mem[16'h1457] = 8'h00;
mem[16'h1458] = 8'h42;
mem[16'h1459] = 8'h22;
mem[16'h145A] = 8'h12;
mem[16'h145B] = 8'h0E;
mem[16'h145C] = 8'h12;
mem[16'h145D] = 8'h22;
mem[16'h145E] = 8'h42;
mem[16'h145F] = 8'h00;
mem[16'h1460] = 8'h02;
mem[16'h1461] = 8'h02;
mem[16'h1462] = 8'h02;
mem[16'h1463] = 8'h02;
mem[16'h1464] = 8'h02;
mem[16'h1465] = 8'h02;
mem[16'h1466] = 8'h7E;
mem[16'h1467] = 8'h00;
mem[16'h1468] = 8'h42;
mem[16'h1469] = 8'h66;
mem[16'h146A] = 8'h5A;
mem[16'h146B] = 8'h5A;
mem[16'h146C] = 8'h42;
mem[16'h146D] = 8'h42;
mem[16'h146E] = 8'h42;
mem[16'h146F] = 8'h00;
mem[16'h1470] = 8'h42;
mem[16'h1471] = 8'h46;
mem[16'h1472] = 8'h4A;
mem[16'h1473] = 8'h52;
mem[16'h1474] = 8'h62;
mem[16'h1475] = 8'h42;
mem[16'h1476] = 8'h42;
mem[16'h1477] = 8'h00;
mem[16'h1478] = 8'h3C;
mem[16'h1479] = 8'h42;
mem[16'h147A] = 8'h42;
mem[16'h147B] = 8'h42;
mem[16'h147C] = 8'h42;
mem[16'h147D] = 8'h42;
mem[16'h147E] = 8'h3C;
mem[16'h147F] = 8'h00;
mem[16'h1480] = 8'h3E;
mem[16'h1481] = 8'h42;
mem[16'h1482] = 8'h42;
mem[16'h1483] = 8'h3E;
mem[16'h1484] = 8'h02;
mem[16'h1485] = 8'h02;
mem[16'h1486] = 8'h02;
mem[16'h1487] = 8'h00;
mem[16'h1488] = 8'h3C;
mem[16'h1489] = 8'h42;
mem[16'h148A] = 8'h42;
mem[16'h148B] = 8'h42;
mem[16'h148C] = 8'h52;
mem[16'h148D] = 8'h22;
mem[16'h148E] = 8'h5C;
mem[16'h148F] = 8'h00;
mem[16'h1490] = 8'h3E;
mem[16'h1491] = 8'h42;
mem[16'h1492] = 8'h42;
mem[16'h1493] = 8'h3E;
mem[16'h1494] = 8'h12;
mem[16'h1495] = 8'h22;
mem[16'h1496] = 8'h42;
mem[16'h1497] = 8'h00;
mem[16'h1498] = 8'h3C;
mem[16'h1499] = 8'h42;
mem[16'h149A] = 8'h02;
mem[16'h149B] = 8'h3C;
mem[16'h149C] = 8'h40;
mem[16'h149D] = 8'h42;
mem[16'h149E] = 8'h3C;
mem[16'h149F] = 8'h00;
mem[16'h14A0] = 8'h7C;
mem[16'h14A1] = 8'h10;
mem[16'h14A2] = 8'h10;
mem[16'h14A3] = 8'h10;
mem[16'h14A4] = 8'h10;
mem[16'h14A5] = 8'h10;
mem[16'h14A6] = 8'h10;
mem[16'h14A7] = 8'h00;
mem[16'h14A8] = 8'h42;
mem[16'h14A9] = 8'h42;
mem[16'h14AA] = 8'h42;
mem[16'h14AB] = 8'h42;
mem[16'h14AC] = 8'h42;
mem[16'h14AD] = 8'h42;
mem[16'h14AE] = 8'h3C;
mem[16'h14AF] = 8'h00;
mem[16'h14B0] = 8'h42;
mem[16'h14B1] = 8'h42;
mem[16'h14B2] = 8'h42;
mem[16'h14B3] = 8'h24;
mem[16'h14B4] = 8'h24;
mem[16'h14B5] = 8'h18;
mem[16'h14B6] = 8'h18;
mem[16'h14B7] = 8'h00;
mem[16'h14B8] = 8'h42;
mem[16'h14B9] = 8'h42;
mem[16'h14BA] = 8'h42;
mem[16'h14BB] = 8'h5A;
mem[16'h14BC] = 8'h5A;
mem[16'h14BD] = 8'h66;
mem[16'h14BE] = 8'h42;
mem[16'h14BF] = 8'h00;
mem[16'h14C0] = 8'h42;
mem[16'h14C1] = 8'h42;
mem[16'h14C2] = 8'h24;
mem[16'h14C3] = 8'h18;
mem[16'h14C4] = 8'h24;
mem[16'h14C5] = 8'h42;
mem[16'h14C6] = 8'h42;
mem[16'h14C7] = 8'h00;
mem[16'h14C8] = 8'h44;
mem[16'h14C9] = 8'h44;
mem[16'h14CA] = 8'h44;
mem[16'h14CB] = 8'h38;
mem[16'h14CC] = 8'h10;
mem[16'h14CD] = 8'h10;
mem[16'h14CE] = 8'h10;
mem[16'h14CF] = 8'h00;
mem[16'h14D0] = 8'h7E;
mem[16'h14D1] = 8'h40;
mem[16'h14D2] = 8'h20;
mem[16'h14D3] = 8'h18;
mem[16'h14D4] = 8'h04;
mem[16'h14D5] = 8'h02;
mem[16'h14D6] = 8'h7E;
mem[16'h14D7] = 8'h00;
mem[16'h14D8] = 8'h3C;
mem[16'h14D9] = 8'h04;
mem[16'h14DA] = 8'h04;
mem[16'h14DB] = 8'h04;
mem[16'h14DC] = 8'h04;
mem[16'h14DD] = 8'h04;
mem[16'h14DE] = 8'h3C;
mem[16'h14DF] = 8'h00;
mem[16'h14E0] = 8'h00;
mem[16'h14E1] = 8'h02;
mem[16'h14E2] = 8'h04;
mem[16'h14E3] = 8'h08;
mem[16'h14E4] = 8'h10;
mem[16'h14E5] = 8'h20;
mem[16'h14E6] = 8'h40;
mem[16'h14E7] = 8'h00;
mem[16'h14E8] = 8'h3C;
mem[16'h14E9] = 8'h20;
mem[16'h14EA] = 8'h20;
mem[16'h14EB] = 8'h20;
mem[16'h14EC] = 8'h20;
mem[16'h14ED] = 8'h20;
mem[16'h14EE] = 8'h3C;
mem[16'h14EF] = 8'h00;
mem[16'h14F0] = 8'h10;
mem[16'h14F1] = 8'h28;
mem[16'h14F2] = 8'h44;
mem[16'h14F3] = 8'h00;
mem[16'h14F4] = 8'h00;
mem[16'h14F5] = 8'h00;
mem[16'h14F6] = 8'h00;
mem[16'h14F7] = 8'h00;
mem[16'h14F8] = 8'h02;
mem[16'h14F9] = 8'h00;
mem[16'h14FA] = 8'h00;
mem[16'h14FB] = 8'h00;
mem[16'h14FC] = 8'h00;
mem[16'h14FD] = 8'h00;
mem[16'h14FE] = 8'h00;
mem[16'h14FF] = 8'hFF;
mem[16'h1500] = 8'h08;
mem[16'h1501] = 8'h10;
mem[16'h1502] = 8'h20;
mem[16'h1503] = 8'h00;
mem[16'h1504] = 8'h00;
mem[16'h1505] = 8'h00;
mem[16'h1506] = 8'h00;
mem[16'h1507] = 8'h00;
mem[16'h1508] = 8'h00;
mem[16'h1509] = 8'h00;
mem[16'h150A] = 8'h1C;
mem[16'h150B] = 8'h20;
mem[16'h150C] = 8'h3C;
mem[16'h150D] = 8'h22;
mem[16'h150E] = 8'h5C;
mem[16'h150F] = 8'h00;
mem[16'h1510] = 8'h02;
mem[16'h1511] = 8'h02;
mem[16'h1512] = 8'h3A;
mem[16'h1513] = 8'h46;
mem[16'h1514] = 8'h42;
mem[16'h1515] = 8'h46;
mem[16'h1516] = 8'h3A;
mem[16'h1517] = 8'h00;
mem[16'h1518] = 8'h00;
mem[16'h1519] = 8'h00;
mem[16'h151A] = 8'h3C;
mem[16'h151B] = 8'h02;
mem[16'h151C] = 8'h02;
mem[16'h151D] = 8'h02;
mem[16'h151E] = 8'h3C;
mem[16'h151F] = 8'h00;
mem[16'h1520] = 8'h40;
mem[16'h1521] = 8'h40;
mem[16'h1522] = 8'h5C;
mem[16'h1523] = 8'h62;
mem[16'h1524] = 8'h42;
mem[16'h1525] = 8'h62;
mem[16'h1526] = 8'h5C;
mem[16'h1527] = 8'h00;
mem[16'h1528] = 8'h00;
mem[16'h1529] = 8'h00;
mem[16'h152A] = 8'h3C;
mem[16'h152B] = 8'h42;
mem[16'h152C] = 8'h7E;
mem[16'h152D] = 8'h02;
mem[16'h152E] = 8'h3C;
mem[16'h152F] = 8'h00;
mem[16'h1530] = 8'h30;
mem[16'h1531] = 8'h48;
mem[16'h1532] = 8'h08;
mem[16'h1533] = 8'h3E;
mem[16'h1534] = 8'h08;
mem[16'h1535] = 8'h08;
mem[16'h1536] = 8'h08;
mem[16'h1537] = 8'h00;
mem[16'h1538] = 8'h00;
mem[16'h1539] = 8'h00;
mem[16'h153A] = 8'h5C;
mem[16'h153B] = 8'h62;
mem[16'h153C] = 8'h62;
mem[16'h153D] = 8'h5C;
mem[16'h153E] = 8'h40;
mem[16'h153F] = 8'h3C;
mem[16'h1540] = 8'h02;
mem[16'h1541] = 8'h02;
mem[16'h1542] = 8'h3A;
mem[16'h1543] = 8'h46;
mem[16'h1544] = 8'h42;
mem[16'h1545] = 8'h42;
mem[16'h1546] = 8'h42;
mem[16'h1547] = 8'h00;
mem[16'h1548] = 8'h10;
mem[16'h1549] = 8'h00;
mem[16'h154A] = 8'h18;
mem[16'h154B] = 8'h10;
mem[16'h154C] = 8'h10;
mem[16'h154D] = 8'h10;
mem[16'h154E] = 8'h38;
mem[16'h154F] = 8'h00;
mem[16'h1550] = 8'h20;
mem[16'h1551] = 8'h00;
mem[16'h1552] = 8'h30;
mem[16'h1553] = 8'h20;
mem[16'h1554] = 8'h20;
mem[16'h1555] = 8'h20;
mem[16'h1556] = 8'h22;
mem[16'h1557] = 8'h1C;
mem[16'h1558] = 8'h02;
mem[16'h1559] = 8'h02;
mem[16'h155A] = 8'h22;
mem[16'h155B] = 8'h12;
mem[16'h155C] = 8'h0A;
mem[16'h155D] = 8'h16;
mem[16'h155E] = 8'h22;
mem[16'h155F] = 8'h00;
mem[16'h1560] = 8'h18;
mem[16'h1561] = 8'h10;
mem[16'h1562] = 8'h10;
mem[16'h1563] = 8'h10;
mem[16'h1564] = 8'h10;
mem[16'h1565] = 8'h10;
mem[16'h1566] = 8'h38;
mem[16'h1567] = 8'h00;
mem[16'h1568] = 8'h00;
mem[16'h1569] = 8'h00;
mem[16'h156A] = 8'h2E;
mem[16'h156B] = 8'h54;
mem[16'h156C] = 8'h54;
mem[16'h156D] = 8'h54;
mem[16'h156E] = 8'h54;
mem[16'h156F] = 8'h00;
mem[16'h1570] = 8'h00;
mem[16'h1571] = 8'h00;
mem[16'h1572] = 8'h3E;
mem[16'h1573] = 8'h44;
mem[16'h1574] = 8'h44;
mem[16'h1575] = 8'h44;
mem[16'h1576] = 8'h44;
mem[16'h1577] = 8'h00;
mem[16'h1578] = 8'h00;
mem[16'h1579] = 8'h00;
mem[16'h157A] = 8'h38;
mem[16'h157B] = 8'h44;
mem[16'h157C] = 8'h44;
mem[16'h157D] = 8'h44;
mem[16'h157E] = 8'h38;
mem[16'h157F] = 8'h00;
mem[16'h1580] = 8'h00;
mem[16'h1581] = 8'h00;
mem[16'h1582] = 8'h3A;
mem[16'h1583] = 8'h46;
mem[16'h1584] = 8'h46;
mem[16'h1585] = 8'h3A;
mem[16'h1586] = 8'h02;
mem[16'h1587] = 8'h02;
mem[16'h1588] = 8'h00;
mem[16'h1589] = 8'h00;
mem[16'h158A] = 8'h5C;
mem[16'h158B] = 8'h62;
mem[16'h158C] = 8'h62;
mem[16'h158D] = 8'h5C;
mem[16'h158E] = 8'h40;
mem[16'h158F] = 8'h40;
mem[16'h1590] = 8'h00;
mem[16'h1591] = 8'h00;
mem[16'h1592] = 8'h3A;
mem[16'h1593] = 8'h46;
mem[16'h1594] = 8'h02;
mem[16'h1595] = 8'h02;
mem[16'h1596] = 8'h02;
mem[16'h1597] = 8'h00;
mem[16'h1598] = 8'h00;
mem[16'h1599] = 8'h00;
mem[16'h159A] = 8'h7C;
mem[16'h159B] = 8'h02;
mem[16'h159C] = 8'h3C;
mem[16'h159D] = 8'h40;
mem[16'h159E] = 8'h3E;
mem[16'h159F] = 8'h00;
mem[16'h15A0] = 8'h08;
mem[16'h15A1] = 8'h08;
mem[16'h15A2] = 8'h3E;
mem[16'h15A3] = 8'h08;
mem[16'h15A4] = 8'h08;
mem[16'h15A5] = 8'h48;
mem[16'h15A6] = 8'h30;
mem[16'h15A7] = 8'h00;
mem[16'h15A8] = 8'h00;
mem[16'h15A9] = 8'h00;
mem[16'h15AA] = 8'h42;
mem[16'h15AB] = 8'h42;
mem[16'h15AC] = 8'h42;
mem[16'h15AD] = 8'h62;
mem[16'h15AE] = 8'h5C;
mem[16'h15AF] = 8'h00;
mem[16'h15B0] = 8'h00;
mem[16'h15B1] = 8'h00;
mem[16'h15B2] = 8'h42;
mem[16'h15B3] = 8'h42;
mem[16'h15B4] = 8'h42;
mem[16'h15B5] = 8'h24;
mem[16'h15B6] = 8'h18;
mem[16'h15B7] = 8'h00;
mem[16'h15B8] = 8'h00;
mem[16'h15B9] = 8'h00;
mem[16'h15BA] = 8'h44;
mem[16'h15BB] = 8'h44;
mem[16'h15BC] = 8'h54;
mem[16'h15BD] = 8'h54;
mem[16'h15BE] = 8'h6C;
mem[16'h15BF] = 8'h00;
mem[16'h15C0] = 8'h00;
mem[16'h15C1] = 8'h00;
mem[16'h15C2] = 8'h42;
mem[16'h15C3] = 8'h24;
mem[16'h15C4] = 8'h18;
mem[16'h15C5] = 8'h24;
mem[16'h15C6] = 8'h42;
mem[16'h15C7] = 8'h00;
mem[16'h15C8] = 8'h00;
mem[16'h15C9] = 8'h00;
mem[16'h15CA] = 8'h42;
mem[16'h15CB] = 8'h42;
mem[16'h15CC] = 8'h62;
mem[16'h15CD] = 8'h5C;
mem[16'h15CE] = 8'h40;
mem[16'h15CF] = 8'h3C;
mem[16'h15D0] = 8'h00;
mem[16'h15D1] = 8'h00;
mem[16'h15D2] = 8'h7E;
mem[16'h15D3] = 8'h20;
mem[16'h15D4] = 8'h18;
mem[16'h15D5] = 8'h04;
mem[16'h15D6] = 8'h7E;
mem[16'h15D7] = 8'h00;
mem[16'h15D8] = 8'h38;
mem[16'h15D9] = 8'h04;
mem[16'h15DA] = 8'h04;
mem[16'h15DB] = 8'h06;
mem[16'h15DC] = 8'h04;
mem[16'h15DD] = 8'h04;
mem[16'h15DE] = 8'h38;
mem[16'h15DF] = 8'h00;
mem[16'h15E0] = 8'h08;
mem[16'h15E1] = 8'h08;
mem[16'h15E2] = 8'h08;
mem[16'h15E3] = 8'h08;
mem[16'h15E4] = 8'h08;
mem[16'h15E5] = 8'h08;
mem[16'h15E6] = 8'h08;
mem[16'h15E7] = 8'h08;
mem[16'h15E8] = 8'h0E;
mem[16'h15E9] = 8'h10;
mem[16'h15EA] = 8'h10;
mem[16'h15EB] = 8'h30;
mem[16'h15EC] = 8'h10;
mem[16'h15ED] = 8'h10;
mem[16'h15EE] = 8'h0E;
mem[16'h15EF] = 8'h00;
mem[16'h15F0] = 8'h28;
mem[16'h15F1] = 8'h14;
mem[16'h15F2] = 8'h00;
mem[16'h15F3] = 8'h00;
mem[16'h15F4] = 8'h00;
mem[16'h15F5] = 8'h00;
mem[16'h15F6] = 8'h00;
mem[16'h15F7] = 8'h00;
mem[16'h15F8] = 8'hFF;
mem[16'h15F9] = 8'hFF;
mem[16'h15FA] = 8'hFF;
mem[16'h15FB] = 8'hFF;
mem[16'h15FC] = 8'hFF;
mem[16'h15FD] = 8'h0F;
mem[16'h15FE] = 8'hAB;
mem[16'h15FF] = 8'h81;
mem[16'h1600] = 8'h30;
mem[16'h1601] = 8'h30;
mem[16'h1602] = 8'h30;
mem[16'h1603] = 8'h30;
mem[16'h1604] = 8'h30;
mem[16'h1605] = 8'h30;
mem[16'h1606] = 8'h30;
mem[16'h1607] = 8'h30;
mem[16'h1608] = 8'h30;
mem[16'h1609] = 8'h30;
mem[16'h160A] = 8'h30;
mem[16'h160B] = 8'h30;
mem[16'h160C] = 8'h30;
mem[16'h160D] = 8'h30;
mem[16'h160E] = 8'h30;
mem[16'h160F] = 8'h30;
mem[16'h1610] = 8'h30;
mem[16'h1611] = 8'h30;
mem[16'h1612] = 8'h30;
mem[16'h1613] = 8'h30;
mem[16'h1614] = 8'h30;
mem[16'h1615] = 8'h30;
mem[16'h1616] = 8'h30;
mem[16'h1617] = 8'h30;
mem[16'h1618] = 8'h30;
mem[16'h1619] = 8'h30;
mem[16'h161A] = 8'h30;
mem[16'h161B] = 8'h30;
mem[16'h161C] = 8'h30;
mem[16'h161D] = 8'h30;
mem[16'h161E] = 8'h30;
mem[16'h161F] = 8'h30;
mem[16'h1620] = 8'h30;
mem[16'h1621] = 8'h30;
mem[16'h1622] = 8'h30;
mem[16'h1623] = 8'h30;
mem[16'h1624] = 8'h30;
mem[16'h1625] = 8'h30;
mem[16'h1626] = 8'h30;
mem[16'h1627] = 8'h30;
mem[16'h1628] = 8'h30;
mem[16'h1629] = 8'h30;
mem[16'h162A] = 8'h30;
mem[16'h162B] = 8'h30;
mem[16'h162C] = 8'h30;
mem[16'h162D] = 8'h30;
mem[16'h162E] = 8'h30;
mem[16'h162F] = 8'h30;
mem[16'h1630] = 8'h30;
mem[16'h1631] = 8'h30;
mem[16'h1632] = 8'h30;
mem[16'h1633] = 8'h30;
mem[16'h1634] = 8'h30;
mem[16'h1635] = 8'h30;
mem[16'h1636] = 8'h30;
mem[16'h1637] = 8'h30;
mem[16'h1638] = 8'h30;
mem[16'h1639] = 8'h30;
mem[16'h163A] = 8'h30;
mem[16'h163B] = 8'h30;
mem[16'h163C] = 8'h30;
mem[16'h163D] = 8'h30;
mem[16'h163E] = 8'h30;
mem[16'h163F] = 8'h30;
mem[16'h1640] = 8'h30;
mem[16'h1641] = 8'h30;
mem[16'h1642] = 8'h30;
mem[16'h1643] = 8'h30;
mem[16'h1644] = 8'h30;
mem[16'h1645] = 8'h30;
mem[16'h1646] = 8'h30;
mem[16'h1647] = 8'h30;
mem[16'h1648] = 8'h30;
mem[16'h1649] = 8'h30;
mem[16'h164A] = 8'h30;
mem[16'h164B] = 8'h30;
mem[16'h164C] = 8'h30;
mem[16'h164D] = 8'h30;
mem[16'h164E] = 8'h30;
mem[16'h164F] = 8'h30;
mem[16'h1650] = 8'h30;
mem[16'h1651] = 8'h30;
mem[16'h1652] = 8'h30;
mem[16'h1653] = 8'h30;
mem[16'h1654] = 8'h30;
mem[16'h1655] = 8'h30;
mem[16'h1656] = 8'h30;
mem[16'h1657] = 8'h30;
mem[16'h1658] = 8'h30;
mem[16'h1659] = 8'h30;
mem[16'h165A] = 8'h30;
mem[16'h165B] = 8'h30;
mem[16'h165C] = 8'h30;
mem[16'h165D] = 8'h30;
mem[16'h165E] = 8'h30;
mem[16'h165F] = 8'h30;
mem[16'h1660] = 8'h30;
mem[16'h1661] = 8'h30;
mem[16'h1662] = 8'h30;
mem[16'h1663] = 8'h30;
mem[16'h1664] = 8'h30;
mem[16'h1665] = 8'h30;
mem[16'h1666] = 8'h30;
mem[16'h1667] = 8'h30;
mem[16'h1668] = 8'h30;
mem[16'h1669] = 8'h30;
mem[16'h166A] = 8'h30;
mem[16'h166B] = 8'h30;
mem[16'h166C] = 8'h30;
mem[16'h166D] = 8'h30;
mem[16'h166E] = 8'h30;
mem[16'h166F] = 8'h30;
mem[16'h1670] = 8'h30;
mem[16'h1671] = 8'h30;
mem[16'h1672] = 8'h30;
mem[16'h1673] = 8'h30;
mem[16'h1674] = 8'h30;
mem[16'h1675] = 8'h30;
mem[16'h1676] = 8'h30;
mem[16'h1677] = 8'h30;
mem[16'h1678] = 8'h30;
mem[16'h1679] = 8'h30;
mem[16'h167A] = 8'h30;
mem[16'h167B] = 8'h30;
mem[16'h167C] = 8'h30;
mem[16'h167D] = 8'h30;
mem[16'h167E] = 8'h30;
mem[16'h167F] = 8'h30;
mem[16'h1680] = 8'h30;
mem[16'h1681] = 8'h30;
mem[16'h1682] = 8'h30;
mem[16'h1683] = 8'h30;
mem[16'h1684] = 8'h30;
mem[16'h1685] = 8'h30;
mem[16'h1686] = 8'h30;
mem[16'h1687] = 8'h30;
mem[16'h1688] = 8'h30;
mem[16'h1689] = 8'h30;
mem[16'h168A] = 8'h30;
mem[16'h168B] = 8'h30;
mem[16'h168C] = 8'h30;
mem[16'h168D] = 8'h30;
mem[16'h168E] = 8'h30;
mem[16'h168F] = 8'h30;
mem[16'h1690] = 8'h30;
mem[16'h1691] = 8'h30;
mem[16'h1692] = 8'h30;
mem[16'h1693] = 8'h30;
mem[16'h1694] = 8'h30;
mem[16'h1695] = 8'h30;
mem[16'h1696] = 8'h30;
mem[16'h1697] = 8'h30;
mem[16'h1698] = 8'h30;
mem[16'h1699] = 8'h30;
mem[16'h169A] = 8'h30;
mem[16'h169B] = 8'h30;
mem[16'h169C] = 8'h30;
mem[16'h169D] = 8'h30;
mem[16'h169E] = 8'h30;
mem[16'h169F] = 8'h30;
mem[16'h16A0] = 8'h30;
mem[16'h16A1] = 8'h30;
mem[16'h16A2] = 8'h30;
mem[16'h16A3] = 8'h30;
mem[16'h16A4] = 8'h30;
mem[16'h16A5] = 8'h30;
mem[16'h16A6] = 8'h30;
mem[16'h16A7] = 8'h30;
mem[16'h16A8] = 8'h30;
mem[16'h16A9] = 8'h30;
mem[16'h16AA] = 8'h30;
mem[16'h16AB] = 8'h30;
mem[16'h16AC] = 8'h30;
mem[16'h16AD] = 8'h30;
mem[16'h16AE] = 8'h30;
mem[16'h16AF] = 8'h30;
mem[16'h16B0] = 8'h30;
mem[16'h16B1] = 8'h30;
mem[16'h16B2] = 8'h30;
mem[16'h16B3] = 8'h30;
mem[16'h16B4] = 8'h30;
mem[16'h16B5] = 8'h30;
mem[16'h16B6] = 8'h30;
mem[16'h16B7] = 8'h30;
mem[16'h16B8] = 8'h30;
mem[16'h16B9] = 8'h30;
mem[16'h16BA] = 8'h30;
mem[16'h16BB] = 8'h30;
mem[16'h16BC] = 8'h30;
mem[16'h16BD] = 8'h30;
mem[16'h16BE] = 8'h30;
mem[16'h16BF] = 8'h30;
mem[16'h16C0] = 8'h30;
mem[16'h16C1] = 8'h30;
mem[16'h16C2] = 8'h30;
mem[16'h16C3] = 8'h30;
mem[16'h16C4] = 8'h30;
mem[16'h16C5] = 8'h30;
mem[16'h16C6] = 8'h30;
mem[16'h16C7] = 8'h30;
mem[16'h16C8] = 8'h30;
mem[16'h16C9] = 8'h30;
mem[16'h16CA] = 8'h30;
mem[16'h16CB] = 8'h30;
mem[16'h16CC] = 8'h30;
mem[16'h16CD] = 8'h30;
mem[16'h16CE] = 8'h30;
mem[16'h16CF] = 8'h30;
mem[16'h16D0] = 8'h30;
mem[16'h16D1] = 8'h30;
mem[16'h16D2] = 8'h30;
mem[16'h16D3] = 8'h30;
mem[16'h16D4] = 8'h30;
mem[16'h16D5] = 8'h30;
mem[16'h16D6] = 8'h30;
mem[16'h16D7] = 8'h30;
mem[16'h16D8] = 8'h30;
mem[16'h16D9] = 8'h30;
mem[16'h16DA] = 8'h30;
mem[16'h16DB] = 8'h30;
mem[16'h16DC] = 8'h30;
mem[16'h16DD] = 8'h30;
mem[16'h16DE] = 8'h30;
mem[16'h16DF] = 8'h30;
mem[16'h16E0] = 8'h30;
mem[16'h16E1] = 8'h30;
mem[16'h16E2] = 8'h30;
mem[16'h16E3] = 8'h30;
mem[16'h16E4] = 8'h30;
mem[16'h16E5] = 8'h30;
mem[16'h16E6] = 8'h30;
mem[16'h16E7] = 8'h30;
mem[16'h16E8] = 8'h30;
mem[16'h16E9] = 8'h30;
mem[16'h16EA] = 8'h30;
mem[16'h16EB] = 8'h30;
mem[16'h16EC] = 8'h30;
mem[16'h16ED] = 8'h30;
mem[16'h16EE] = 8'h30;
mem[16'h16EF] = 8'h30;
mem[16'h16F0] = 8'h30;
mem[16'h16F1] = 8'h30;
mem[16'h16F2] = 8'h30;
mem[16'h16F3] = 8'h30;
mem[16'h16F4] = 8'h30;
mem[16'h16F5] = 8'h30;
mem[16'h16F6] = 8'h30;
mem[16'h16F7] = 8'h30;
mem[16'h16F8] = 8'h30;
mem[16'h16F9] = 8'h30;
mem[16'h16FA] = 8'h30;
mem[16'h16FB] = 8'h30;
mem[16'h16FC] = 8'h30;
mem[16'h16FD] = 8'h00;
mem[16'h16FE] = 8'h00;
mem[16'h16FF] = 8'h00;
mem[16'h1700] = 8'hA0;
mem[16'h1701] = 8'h03;
mem[16'h1702] = 8'h84;
mem[16'h1703] = 8'h37;
mem[16'h1704] = 8'hA0;
mem[16'h1705] = 8'h09;
mem[16'h1706] = 8'h84;
mem[16'h1707] = 8'h36;
mem[16'h1708] = 8'h60;
mem[16'h1709] = 8'h48;
mem[16'h170A] = 8'h84;
mem[16'h170B] = 8'h4E;
mem[16'h170C] = 8'hC9;
mem[16'h170D] = 8'h8D;
mem[16'h170E] = 8'hF0;
mem[16'h170F] = 8'h68;
mem[16'h1710] = 8'hA5;
mem[16'h1711] = 8'h25;
mem[16'h1712] = 8'h4A;
mem[16'h1713] = 8'h29;
mem[16'h1714] = 8'h03;
mem[16'h1715] = 8'h09;
mem[16'h1716] = 8'h20;
mem[16'h1717] = 8'h85;
mem[16'h1718] = 8'h2B;
mem[16'h1719] = 8'hA5;
mem[16'h171A] = 8'h25;
mem[16'h171B] = 8'h6A;
mem[16'h171C] = 8'h08;
mem[16'h171D] = 8'h0A;
mem[16'h171E] = 8'h29;
mem[16'h171F] = 8'h18;
mem[16'h1720] = 8'h85;
mem[16'h1721] = 8'h2A;
mem[16'h1722] = 8'h0A;
mem[16'h1723] = 8'h0A;
mem[16'h1724] = 8'h05;
mem[16'h1725] = 8'h2A;
mem[16'h1726] = 8'h0A;
mem[16'h1727] = 8'h28;
mem[16'h1728] = 8'h6A;
mem[16'h1729] = 8'h18;
mem[16'h172A] = 8'h65;
mem[16'h172B] = 8'h24;
mem[16'h172C] = 8'h85;
mem[16'h172D] = 8'h2A;
mem[16'h172E] = 8'h68;
mem[16'h172F] = 8'h29;
mem[16'h1730] = 8'h7F;
mem[16'h1731] = 8'h48;
mem[16'h1732] = 8'hA9;
mem[16'h1733] = 8'h00;
mem[16'h1734] = 8'h85;
mem[16'h1735] = 8'h27;
mem[16'h1736] = 8'h68;
mem[16'h1737] = 8'h48;
mem[16'h1738] = 8'h2A;
mem[16'h1739] = 8'h26;
mem[16'h173A] = 8'h27;
mem[16'h173B] = 8'h2A;
mem[16'h173C] = 8'h26;
mem[16'h173D] = 8'h27;
mem[16'h173E] = 8'h2A;
mem[16'h173F] = 8'h26;
mem[16'h1740] = 8'h27;
mem[16'h1741] = 8'h85;
mem[16'h1742] = 8'h26;
mem[16'h1743] = 8'hA5;
mem[16'h1744] = 8'h27;
mem[16'h1745] = 8'h18;
mem[16'h1746] = 8'h69;
mem[16'h1747] = 8'h04;
mem[16'h1748] = 8'h85;
mem[16'h1749] = 8'h27;
mem[16'h174A] = 8'hA0;
mem[16'h174B] = 8'h00;
mem[16'h174C] = 8'hB1;
mem[16'h174D] = 8'h26;
mem[16'h174E] = 8'h48;
mem[16'h174F] = 8'h84;
mem[16'h1750] = 8'h4F;
mem[16'h1751] = 8'hA0;
mem[16'h1752] = 8'h00;
mem[16'h1753] = 8'h51;
mem[16'h1754] = 8'h2A;
mem[16'h1755] = 8'h91;
mem[16'h1756] = 8'h2A;
mem[16'h1757] = 8'hA5;
mem[16'h1758] = 8'h2B;
mem[16'h1759] = 8'hEA;
mem[16'h175A] = 8'hEA;
mem[16'h175B] = 8'h85;
mem[16'h175C] = 8'h2B;
mem[16'h175D] = 8'h68;
mem[16'h175E] = 8'h51;
mem[16'h175F] = 8'h2A;
mem[16'h1760] = 8'hEA;
mem[16'h1761] = 8'hEA;
mem[16'h1762] = 8'hA4;
mem[16'h1763] = 8'h4F;
mem[16'h1764] = 8'hA5;
mem[16'h1765] = 8'h2B;
mem[16'h1766] = 8'h18;
mem[16'h1767] = 8'h69;
mem[16'h1768] = 8'h04;
mem[16'h1769] = 8'h85;
mem[16'h176A] = 8'h2B;
mem[16'h176B] = 8'hC8;
mem[16'h176C] = 8'hC0;
mem[16'h176D] = 8'h08;
mem[16'h176E] = 8'hD0;
mem[16'h176F] = 8'hDC;
mem[16'h1770] = 8'hE6;
mem[16'h1771] = 8'h24;
mem[16'h1772] = 8'hA5;
mem[16'h1773] = 8'h24;
mem[16'h1774] = 8'hC5;
mem[16'h1775] = 8'h21;
mem[16'h1776] = 8'h90;
mem[16'h1777] = 8'h10;
mem[16'h1778] = 8'hA5;
mem[16'h1779] = 8'h20;
mem[16'h177A] = 8'h85;
mem[16'h177B] = 8'h24;
mem[16'h177C] = 8'hE6;
mem[16'h177D] = 8'h25;
mem[16'h177E] = 8'hA5;
mem[16'h177F] = 8'h25;
mem[16'h1780] = 8'hC5;
mem[16'h1781] = 8'h23;
mem[16'h1782] = 8'h90;
mem[16'h1783] = 8'h04;
mem[16'h1784] = 8'hA5;
mem[16'h1785] = 8'h22;
mem[16'h1786] = 8'h85;
mem[16'h1787] = 8'h25;
mem[16'h1788] = 8'hA4;
mem[16'h1789] = 8'h4E;
mem[16'h178A] = 8'h68;
mem[16'h178B] = 8'h60;
mem[16'h178C] = 8'hFF;
mem[16'h178D] = 8'hFF;
mem[16'h178E] = 8'h00;
mem[16'h178F] = 8'h00;
mem[16'h1790] = 8'hFF;
mem[16'h1791] = 8'hFF;
mem[16'h1792] = 8'h00;
mem[16'h1793] = 8'h00;
mem[16'h1794] = 8'hFF;
mem[16'h1795] = 8'hFF;
mem[16'h1796] = 8'h00;
mem[16'h1797] = 8'h00;
mem[16'h1798] = 8'hFF;
mem[16'h1799] = 8'hFF;
mem[16'h179A] = 8'h00;
mem[16'h179B] = 8'h00;
mem[16'h179C] = 8'hFF;
mem[16'h179D] = 8'hFF;
mem[16'h179E] = 8'h00;
mem[16'h179F] = 8'h00;
mem[16'h17A0] = 8'hFF;
mem[16'h17A1] = 8'hFF;
mem[16'h17A2] = 8'h00;
mem[16'h17A3] = 8'h00;
mem[16'h17A4] = 8'hFF;
mem[16'h17A5] = 8'hFF;
mem[16'h17A6] = 8'h00;
mem[16'h17A7] = 8'h00;
mem[16'h17A8] = 8'hFF;
mem[16'h17A9] = 8'hFF;
mem[16'h17AA] = 8'h00;
mem[16'h17AB] = 8'h00;
mem[16'h17AC] = 8'hFF;
mem[16'h17AD] = 8'hFF;
mem[16'h17AE] = 8'h00;
mem[16'h17AF] = 8'h00;
mem[16'h17B0] = 8'hFF;
mem[16'h17B1] = 8'hFF;
mem[16'h17B2] = 8'h00;
mem[16'h17B3] = 8'h00;
mem[16'h17B4] = 8'hFF;
mem[16'h17B5] = 8'hFF;
mem[16'h17B6] = 8'h00;
mem[16'h17B7] = 8'h00;
mem[16'h17B8] = 8'hFF;
mem[16'h17B9] = 8'hFF;
mem[16'h17BA] = 8'h00;
mem[16'h17BB] = 8'h00;
mem[16'h17BC] = 8'hFF;
mem[16'h17BD] = 8'hFF;
mem[16'h17BE] = 8'h00;
mem[16'h17BF] = 8'h00;
mem[16'h17C0] = 8'h00;
mem[16'h17C1] = 8'h00;
mem[16'h17C2] = 8'h00;
mem[16'h17C3] = 8'h00;
mem[16'h17C4] = 8'h00;
mem[16'h17C5] = 8'h00;
mem[16'h17C6] = 8'h00;
mem[16'h17C7] = 8'h00;
mem[16'h17C8] = 8'h00;
mem[16'h17C9] = 8'h00;
mem[16'h17CA] = 8'h00;
mem[16'h17CB] = 8'h00;
mem[16'h17CC] = 8'hB6;
mem[16'h17CD] = 8'h00;
mem[16'h17CE] = 8'h00;
mem[16'h17CF] = 8'h00;
mem[16'h17D0] = 8'h4C;
mem[16'h17D1] = 8'hBF;
mem[16'h17D2] = 8'h9D;
mem[16'h17D3] = 8'h4C;
mem[16'h17D4] = 8'h84;
mem[16'h17D5] = 8'h9D;
mem[16'h17D6] = 8'h4C;
mem[16'h17D7] = 8'hFD;
mem[16'h17D8] = 8'hAA;
mem[16'h17D9] = 8'h4C;
mem[16'h17DA] = 8'hB5;
mem[16'h17DB] = 8'hB7;
mem[16'h17DC] = 8'hAD;
mem[16'h17DD] = 8'h0F;
mem[16'h17DE] = 8'h9D;
mem[16'h17DF] = 8'hAC;
mem[16'h17E0] = 8'h0E;
mem[16'h17E1] = 8'h9D;
mem[16'h17E2] = 8'h60;
mem[16'h17E3] = 8'hAD;
mem[16'h17E4] = 8'hC2;
mem[16'h17E5] = 8'hAA;
mem[16'h17E6] = 8'hAC;
mem[16'h17E7] = 8'hC1;
mem[16'h17E8] = 8'hAA;
mem[16'h17E9] = 8'h60;
mem[16'h17EA] = 8'h4C;
mem[16'h17EB] = 8'h51;
mem[16'h17EC] = 8'hA8;
mem[16'h17ED] = 8'hEA;
mem[16'h17EE] = 8'hEA;
mem[16'h17EF] = 8'h4C;
mem[16'h17F0] = 8'h59;
mem[16'h17F1] = 8'hFA;
mem[16'h17F2] = 8'h43;
mem[16'h17F3] = 8'h30;
mem[16'h17F4] = 8'h95;
mem[16'h17F5] = 8'h4C;
mem[16'h17F6] = 8'h58;
mem[16'h17F7] = 8'hFF;
mem[16'h17F8] = 8'h4C;
mem[16'h17F9] = 8'h65;
mem[16'h17FA] = 8'hFF;
mem[16'h17FB] = 8'h4C;
mem[16'h17FC] = 8'h65;
mem[16'h17FD] = 8'hFF;
mem[16'h17FE] = 8'h65;
mem[16'h17FF] = 8'hFF;
mem[16'h1800] = 8'h00;
mem[16'h1801] = 8'hFF;
mem[16'h1802] = 8'hFF;
mem[16'h1803] = 8'h00;
mem[16'h1804] = 8'h00;
mem[16'h1805] = 8'hFF;
mem[16'h1806] = 8'hFF;
mem[16'h1807] = 8'h00;
mem[16'h1808] = 8'h00;
mem[16'h1809] = 8'hFF;
mem[16'h180A] = 8'hFF;
mem[16'h180B] = 8'h00;
mem[16'h180C] = 8'h00;
mem[16'h180D] = 8'hFF;
mem[16'h180E] = 8'hFF;
mem[16'h180F] = 8'h00;
mem[16'h1810] = 8'h00;
mem[16'h1811] = 8'hFF;
mem[16'h1812] = 8'hFF;
mem[16'h1813] = 8'h00;
mem[16'h1814] = 8'h00;
mem[16'h1815] = 8'hFF;
mem[16'h1816] = 8'hFF;
mem[16'h1817] = 8'h00;
mem[16'h1818] = 8'h00;
mem[16'h1819] = 8'hFF;
mem[16'h181A] = 8'hFF;
mem[16'h181B] = 8'h00;
mem[16'h181C] = 8'h00;
mem[16'h181D] = 8'hFF;
mem[16'h181E] = 8'hFF;
mem[16'h181F] = 8'h00;
mem[16'h1820] = 8'h00;
mem[16'h1821] = 8'hFF;
mem[16'h1822] = 8'hFF;
mem[16'h1823] = 8'h00;
mem[16'h1824] = 8'h00;
mem[16'h1825] = 8'hFF;
mem[16'h1826] = 8'hFF;
mem[16'h1827] = 8'h00;
mem[16'h1828] = 8'h00;
mem[16'h1829] = 8'hFF;
mem[16'h182A] = 8'hFF;
mem[16'h182B] = 8'h00;
mem[16'h182C] = 8'h00;
mem[16'h182D] = 8'hFF;
mem[16'h182E] = 8'hFF;
mem[16'h182F] = 8'h00;
mem[16'h1830] = 8'h00;
mem[16'h1831] = 8'hFF;
mem[16'h1832] = 8'hFF;
mem[16'h1833] = 8'h00;
mem[16'h1834] = 8'h00;
mem[16'h1835] = 8'hFF;
mem[16'h1836] = 8'hFF;
mem[16'h1837] = 8'h00;
mem[16'h1838] = 8'h00;
mem[16'h1839] = 8'h14;
mem[16'h183A] = 8'h22;
mem[16'h183B] = 8'h22;
mem[16'h183C] = 8'h22;
mem[16'h183D] = 8'h41;
mem[16'h183E] = 8'h7F;
mem[16'h183F] = 8'h08;
mem[16'h1840] = 8'h10;
mem[16'h1841] = 8'h08;
mem[16'h1842] = 8'h04;
mem[16'h1843] = 8'h7E;
mem[16'h1844] = 8'h04;
mem[16'h1845] = 8'h08;
mem[16'h1846] = 8'h10;
mem[16'h1847] = 8'h00;
mem[16'h1848] = 8'h08;
mem[16'h1849] = 8'h10;
mem[16'h184A] = 8'h20;
mem[16'h184B] = 8'h7E;
mem[16'h184C] = 8'h20;
mem[16'h184D] = 8'h10;
mem[16'h184E] = 8'h08;
mem[16'h184F] = 8'h00;
mem[16'h1850] = 8'h08;
mem[16'h1851] = 8'h08;
mem[16'h1852] = 8'h08;
mem[16'h1853] = 8'h49;
mem[16'h1854] = 8'h2A;
mem[16'h1855] = 8'h1C;
mem[16'h1856] = 8'h08;
mem[16'h1857] = 8'h00;
mem[16'h1858] = 8'h08;
mem[16'h1859] = 8'h1C;
mem[16'h185A] = 8'h2A;
mem[16'h185B] = 8'h49;
mem[16'h185C] = 8'h08;
mem[16'h185D] = 8'h08;
mem[16'h185E] = 8'h08;
mem[16'h185F] = 8'h00;
mem[16'h1860] = 8'h08;
mem[16'h1861] = 8'h49;
mem[16'h1862] = 8'h2A;
mem[16'h1863] = 8'h1C;
mem[16'h1864] = 8'h49;
mem[16'h1865] = 8'h2A;
mem[16'h1866] = 8'h1C;
mem[16'h1867] = 8'h08;
mem[16'h1868] = 8'h40;
mem[16'h1869] = 8'h60;
mem[16'h186A] = 8'h70;
mem[16'h186B] = 8'h78;
mem[16'h186C] = 8'h70;
mem[16'h186D] = 8'h60;
mem[16'h186E] = 8'h40;
mem[16'h186F] = 8'h00;
mem[16'h1870] = 8'h40;
mem[16'h1871] = 8'h40;
mem[16'h1872] = 8'h20;
mem[16'h1873] = 8'h20;
mem[16'h1874] = 8'h13;
mem[16'h1875] = 8'h14;
mem[16'h1876] = 8'h0C;
mem[16'h1877] = 8'h08;
mem[16'h1878] = 8'h1A;
mem[16'h1879] = 8'h00;
mem[16'h187A] = 8'h00;
mem[16'h187B] = 8'h7C;
mem[16'h187C] = 8'h2A;
mem[16'h187D] = 8'h28;
mem[16'h187E] = 8'h34;
mem[16'h187F] = 8'h00;
mem[16'h1880] = 8'h36;
mem[16'h1881] = 8'h7F;
mem[16'h1882] = 8'h7F;
mem[16'h1883] = 8'h7F;
mem[16'h1884] = 8'h3E;
mem[16'h1885] = 8'h1C;
mem[16'h1886] = 8'h08;
mem[16'h1887] = 8'h00;
mem[16'h1888] = 8'h08;
mem[16'h1889] = 8'h1C;
mem[16'h188A] = 8'h3E;
mem[16'h188B] = 8'h7F;
mem[16'h188C] = 8'h3E;
mem[16'h188D] = 8'h1C;
mem[16'h188E] = 8'h08;
mem[16'h188F] = 8'h00;
mem[16'h1890] = 8'h08;
mem[16'h1891] = 8'h1C;
mem[16'h1892] = 8'h3E;
mem[16'h1893] = 8'h7F;
mem[16'h1894] = 8'h7F;
mem[16'h1895] = 8'h2A;
mem[16'h1896] = 8'h08;
mem[16'h1897] = 8'h00;
mem[16'h1898] = 8'h08;
mem[16'h1899] = 8'h1C;
mem[16'h189A] = 8'h1C;
mem[16'h189B] = 8'h2A;
mem[16'h189C] = 8'h7F;
mem[16'h189D] = 8'h7F;
mem[16'h189E] = 8'h2A;
mem[16'h189F] = 8'h08;
mem[16'h18A0] = 8'h3E;
mem[16'h18A1] = 8'h08;
mem[16'h18A2] = 8'h08;
mem[16'h18A3] = 8'h22;
mem[16'h18A4] = 8'h36;
mem[16'h18A5] = 8'h2A;
mem[16'h18A6] = 8'h22;
mem[16'h18A7] = 8'h00;
mem[16'h18A8] = 8'h00;
mem[16'h18A9] = 8'h22;
mem[16'h18AA] = 8'h14;
mem[16'h18AB] = 8'h08;
mem[16'h18AC] = 8'h14;
mem[16'h18AD] = 8'h22;
mem[16'h18AE] = 8'h00;
mem[16'h18AF] = 8'h00;
mem[16'h18B0] = 8'h04;
mem[16'h18B1] = 8'h0E;
mem[16'h18B2] = 8'h04;
mem[16'h18B3] = 8'h04;
mem[16'h18B4] = 8'h00;
mem[16'h18B5] = 8'h00;
mem[16'h18B6] = 8'h00;
mem[16'h18B7] = 8'h00;
mem[16'h18B8] = 8'h00;
mem[16'h18B9] = 8'h08;
mem[16'h18BA] = 8'h00;
mem[16'h18BB] = 8'h3E;
mem[16'h18BC] = 8'h00;
mem[16'h18BD] = 8'h08;
mem[16'h18BE] = 8'h00;
mem[16'h18BF] = 8'h00;
mem[16'h18C0] = 8'h18;
mem[16'h18C1] = 8'h24;
mem[16'h18C2] = 8'h08;
mem[16'h18C3] = 8'h14;
mem[16'h18C4] = 8'h08;
mem[16'h18C5] = 8'h12;
mem[16'h18C6] = 8'h0C;
mem[16'h18C7] = 8'h00;
mem[16'h18C8] = 8'h10;
mem[16'h18C9] = 8'h38;
mem[16'h18CA] = 8'h04;
mem[16'h18CB] = 8'h04;
mem[16'h18CC] = 8'h38;
mem[16'h18CD] = 8'h10;
mem[16'h18CE] = 8'h00;
mem[16'h18CF] = 8'h00;
mem[16'h18D0] = 8'h08;
mem[16'h18D1] = 8'h1C;
mem[16'h18D2] = 8'h08;
mem[16'h18D3] = 8'h1C;
mem[16'h18D4] = 8'h3E;
mem[16'h18D5] = 8'h1C;
mem[16'h18D6] = 8'h3E;
mem[16'h18D7] = 8'h7F;
mem[16'h18D8] = 8'h08;
mem[16'h18D9] = 8'h3E;
mem[16'h18DA] = 8'h1C;
mem[16'h18DB] = 8'h08;
mem[16'h18DC] = 8'h1C;
mem[16'h18DD] = 8'h1C;
mem[16'h18DE] = 8'h3E;
mem[16'h18DF] = 8'h7F;
mem[16'h18E0] = 8'h00;
mem[16'h18E1] = 8'h2A;
mem[16'h18E2] = 8'h3E;
mem[16'h18E3] = 8'h1C;
mem[16'h18E4] = 8'h1C;
mem[16'h18E5] = 8'h1C;
mem[16'h18E6] = 8'h3E;
mem[16'h18E7] = 8'h7F;
mem[16'h18E8] = 8'h00;
mem[16'h18E9] = 8'h10;
mem[16'h18EA] = 8'h3C;
mem[16'h18EB] = 8'h3E;
mem[16'h18EC] = 8'h18;
mem[16'h18ED] = 8'h0C;
mem[16'h18EE] = 8'h1E;
mem[16'h18EF] = 8'h3F;
mem[16'h18F0] = 8'h00;
mem[16'h18F1] = 8'h08;
mem[16'h18F2] = 8'h18;
mem[16'h18F3] = 8'h3A;
mem[16'h18F4] = 8'h7B;
mem[16'h18F5] = 8'h3E;
mem[16'h18F6] = 8'h1C;
mem[16'h18F7] = 8'h7F;
mem[16'h18F8] = 8'h04;
mem[16'h18F9] = 8'h00;
mem[16'h18FA] = 8'h08;
mem[16'h18FB] = 8'h1C;
mem[16'h18FC] = 8'h1C;
mem[16'h18FD] = 8'h08;
mem[16'h18FE] = 8'h1C;
mem[16'h18FF] = 8'h3E;
mem[16'h1900] = 8'h00;
mem[16'h1901] = 8'h00;
mem[16'h1902] = 8'h00;
mem[16'h1903] = 8'h00;
mem[16'h1904] = 8'h00;
mem[16'h1905] = 8'h00;
mem[16'h1906] = 8'h00;
mem[16'h1907] = 8'h00;
mem[16'h1908] = 8'h10;
mem[16'h1909] = 8'h10;
mem[16'h190A] = 8'h10;
mem[16'h190B] = 8'h10;
mem[16'h190C] = 8'h00;
mem[16'h190D] = 8'h00;
mem[16'h190E] = 8'h10;
mem[16'h190F] = 8'h00;
mem[16'h1910] = 8'h24;
mem[16'h1911] = 8'h24;
mem[16'h1912] = 8'h24;
mem[16'h1913] = 8'h00;
mem[16'h1914] = 8'h00;
mem[16'h1915] = 8'h00;
mem[16'h1916] = 8'h00;
mem[16'h1917] = 8'h00;
mem[16'h1918] = 8'h24;
mem[16'h1919] = 8'h24;
mem[16'h191A] = 8'h7E;
mem[16'h191B] = 8'h24;
mem[16'h191C] = 8'h7E;
mem[16'h191D] = 8'h24;
mem[16'h191E] = 8'h24;
mem[16'h191F] = 8'h00;
mem[16'h1920] = 8'h10;
mem[16'h1921] = 8'h78;
mem[16'h1922] = 8'h14;
mem[16'h1923] = 8'h38;
mem[16'h1924] = 8'h50;
mem[16'h1925] = 8'h3C;
mem[16'h1926] = 8'h10;
mem[16'h1927] = 8'h00;
mem[16'h1928] = 8'h00;
mem[16'h1929] = 8'h46;
mem[16'h192A] = 8'h26;
mem[16'h192B] = 8'h10;
mem[16'h192C] = 8'h08;
mem[16'h192D] = 8'h64;
mem[16'h192E] = 8'h62;
mem[16'h192F] = 8'h00;
mem[16'h1930] = 8'h0C;
mem[16'h1931] = 8'h12;
mem[16'h1932] = 8'h12;
mem[16'h1933] = 8'h0C;
mem[16'h1934] = 8'h52;
mem[16'h1935] = 8'h22;
mem[16'h1936] = 8'h5C;
mem[16'h1937] = 8'h00;
mem[16'h1938] = 8'h20;
mem[16'h1939] = 8'h10;
mem[16'h193A] = 8'h08;
mem[16'h193B] = 8'h00;
mem[16'h193C] = 8'h00;
mem[16'h193D] = 8'h00;
mem[16'h193E] = 8'h00;
mem[16'h193F] = 8'h00;
mem[16'h1940] = 8'h20;
mem[16'h1941] = 8'h10;
mem[16'h1942] = 8'h08;
mem[16'h1943] = 8'h08;
mem[16'h1944] = 8'h08;
mem[16'h1945] = 8'h10;
mem[16'h1946] = 8'h20;
mem[16'h1947] = 8'h00;
mem[16'h1948] = 8'h04;
mem[16'h1949] = 8'h08;
mem[16'h194A] = 8'h10;
mem[16'h194B] = 8'h10;
mem[16'h194C] = 8'h10;
mem[16'h194D] = 8'h08;
mem[16'h194E] = 8'h04;
mem[16'h194F] = 8'h00;
mem[16'h1950] = 8'h10;
mem[16'h1951] = 8'h54;
mem[16'h1952] = 8'h38;
mem[16'h1953] = 8'h7C;
mem[16'h1954] = 8'h38;
mem[16'h1955] = 8'h54;
mem[16'h1956] = 8'h10;
mem[16'h1957] = 8'h00;
mem[16'h1958] = 8'h00;
mem[16'h1959] = 8'h10;
mem[16'h195A] = 8'h10;
mem[16'h195B] = 8'h7C;
mem[16'h195C] = 8'h10;
mem[16'h195D] = 8'h10;
mem[16'h195E] = 8'h00;
mem[16'h195F] = 8'h00;
mem[16'h1960] = 8'h00;
mem[16'h1961] = 8'h00;
mem[16'h1962] = 8'h00;
mem[16'h1963] = 8'h00;
mem[16'h1964] = 8'h00;
mem[16'h1965] = 8'h18;
mem[16'h1966] = 8'h18;
mem[16'h1967] = 8'h0C;
mem[16'h1968] = 8'h00;
mem[16'h1969] = 8'h00;
mem[16'h196A] = 8'h00;
mem[16'h196B] = 8'h7E;
mem[16'h196C] = 8'h00;
mem[16'h196D] = 8'h00;
mem[16'h196E] = 8'h00;
mem[16'h196F] = 8'h00;
mem[16'h1970] = 8'h00;
mem[16'h1971] = 8'h00;
mem[16'h1972] = 8'h00;
mem[16'h1973] = 8'h00;
mem[16'h1974] = 8'h00;
mem[16'h1975] = 8'h18;
mem[16'h1976] = 8'h18;
mem[16'h1977] = 8'h00;
mem[16'h1978] = 8'h28;
mem[16'h1979] = 8'h40;
mem[16'h197A] = 8'h20;
mem[16'h197B] = 8'h10;
mem[16'h197C] = 8'h08;
mem[16'h197D] = 8'h04;
mem[16'h197E] = 8'h02;
mem[16'h197F] = 8'h00;
mem[16'h1980] = 8'h3C;
mem[16'h1981] = 8'h42;
mem[16'h1982] = 8'h42;
mem[16'h1983] = 8'h42;
mem[16'h1984] = 8'h42;
mem[16'h1985] = 8'h42;
mem[16'h1986] = 8'h3C;
mem[16'h1987] = 8'h00;
mem[16'h1988] = 8'h10;
mem[16'h1989] = 8'h18;
mem[16'h198A] = 8'h14;
mem[16'h198B] = 8'h10;
mem[16'h198C] = 8'h10;
mem[16'h198D] = 8'h10;
mem[16'h198E] = 8'h7C;
mem[16'h198F] = 8'h00;
mem[16'h1990] = 8'h3C;
mem[16'h1991] = 8'h42;
mem[16'h1992] = 8'h40;
mem[16'h1993] = 8'h30;
mem[16'h1994] = 8'h0C;
mem[16'h1995] = 8'h02;
mem[16'h1996] = 8'h7E;
mem[16'h1997] = 8'h00;
mem[16'h1998] = 8'h3C;
mem[16'h1999] = 8'h42;
mem[16'h199A] = 8'h40;
mem[16'h199B] = 8'h38;
mem[16'h199C] = 8'h40;
mem[16'h199D] = 8'h42;
mem[16'h199E] = 8'h3C;
mem[16'h199F] = 8'h00;
mem[16'h19A0] = 8'h20;
mem[16'h19A1] = 8'h30;
mem[16'h19A2] = 8'h28;
mem[16'h19A3] = 8'h24;
mem[16'h19A4] = 8'h7E;
mem[16'h19A5] = 8'h20;
mem[16'h19A6] = 8'h20;
mem[16'h19A7] = 8'h00;
mem[16'h19A8] = 8'h7E;
mem[16'h19A9] = 8'h02;
mem[16'h19AA] = 8'h1E;
mem[16'h19AB] = 8'h20;
mem[16'h19AC] = 8'h40;
mem[16'h19AD] = 8'h22;
mem[16'h19AE] = 8'h1C;
mem[16'h19AF] = 8'h00;
mem[16'h19B0] = 8'h38;
mem[16'h19B1] = 8'h04;
mem[16'h19B2] = 8'h02;
mem[16'h19B3] = 8'h3E;
mem[16'h19B4] = 8'h42;
mem[16'h19B5] = 8'h42;
mem[16'h19B6] = 8'h3C;
mem[16'h19B7] = 8'h00;
mem[16'h19B8] = 8'h7E;
mem[16'h19B9] = 8'h42;
mem[16'h19BA] = 8'h20;
mem[16'h19BB] = 8'h10;
mem[16'h19BC] = 8'h08;
mem[16'h19BD] = 8'h08;
mem[16'h19BE] = 8'h08;
mem[16'h19BF] = 8'h00;
mem[16'h19C0] = 8'h3C;
mem[16'h19C1] = 8'h42;
mem[16'h19C2] = 8'h42;
mem[16'h19C3] = 8'h3C;
mem[16'h19C4] = 8'h42;
mem[16'h19C5] = 8'h42;
mem[16'h19C6] = 8'h3C;
mem[16'h19C7] = 8'h00;
mem[16'h19C8] = 8'h3C;
mem[16'h19C9] = 8'h42;
mem[16'h19CA] = 8'h42;
mem[16'h19CB] = 8'h7C;
mem[16'h19CC] = 8'h40;
mem[16'h19CD] = 8'h20;
mem[16'h19CE] = 8'h1C;
mem[16'h19CF] = 8'h00;
mem[16'h19D0] = 8'h00;
mem[16'h19D1] = 8'h00;
mem[16'h19D2] = 8'h18;
mem[16'h19D3] = 8'h18;
mem[16'h19D4] = 8'h00;
mem[16'h19D5] = 8'h18;
mem[16'h19D6] = 8'h18;
mem[16'h19D7] = 8'h00;
mem[16'h19D8] = 8'h00;
mem[16'h19D9] = 8'h00;
mem[16'h19DA] = 8'h18;
mem[16'h19DB] = 8'h18;
mem[16'h19DC] = 8'h00;
mem[16'h19DD] = 8'h18;
mem[16'h19DE] = 8'h18;
mem[16'h19DF] = 8'h0C;
mem[16'h19E0] = 8'h20;
mem[16'h19E1] = 8'h10;
mem[16'h19E2] = 8'h08;
mem[16'h19E3] = 8'h04;
mem[16'h19E4] = 8'h08;
mem[16'h19E5] = 8'h10;
mem[16'h19E6] = 8'h20;
mem[16'h19E7] = 8'h00;
mem[16'h19E8] = 8'h00;
mem[16'h19E9] = 8'h00;
mem[16'h19EA] = 8'h3E;
mem[16'h19EB] = 8'h00;
mem[16'h19EC] = 8'h3E;
mem[16'h19ED] = 8'h00;
mem[16'h19EE] = 8'h00;
mem[16'h19EF] = 8'h00;
mem[16'h19F0] = 8'h04;
mem[16'h19F1] = 8'h08;
mem[16'h19F2] = 8'h10;
mem[16'h19F3] = 8'h20;
mem[16'h19F4] = 8'h10;
mem[16'h19F5] = 8'h08;
mem[16'h19F6] = 8'h04;
mem[16'h19F7] = 8'h00;
mem[16'h19F8] = 8'h60;
mem[16'h19F9] = 8'h42;
mem[16'h19FA] = 8'h40;
mem[16'h19FB] = 8'h30;
mem[16'h19FC] = 8'h08;
mem[16'h19FD] = 8'h00;
mem[16'h19FE] = 8'h08;
mem[16'h19FF] = 8'h00;
mem[16'h1A00] = 8'h38;
mem[16'h1A01] = 8'h44;
mem[16'h1A02] = 8'h52;
mem[16'h1A03] = 8'h6A;
mem[16'h1A04] = 8'h32;
mem[16'h1A05] = 8'h04;
mem[16'h1A06] = 8'h78;
mem[16'h1A07] = 8'h00;
mem[16'h1A08] = 8'h18;
mem[16'h1A09] = 8'h24;
mem[16'h1A0A] = 8'h42;
mem[16'h1A0B] = 8'h7E;
mem[16'h1A0C] = 8'h42;
mem[16'h1A0D] = 8'h42;
mem[16'h1A0E] = 8'h42;
mem[16'h1A0F] = 8'h00;
mem[16'h1A10] = 8'h3E;
mem[16'h1A11] = 8'h44;
mem[16'h1A12] = 8'h44;
mem[16'h1A13] = 8'h3C;
mem[16'h1A14] = 8'h44;
mem[16'h1A15] = 8'h44;
mem[16'h1A16] = 8'h3E;
mem[16'h1A17] = 8'h00;
mem[16'h1A18] = 8'h3C;
mem[16'h1A19] = 8'h42;
mem[16'h1A1A] = 8'h02;
mem[16'h1A1B] = 8'h02;
mem[16'h1A1C] = 8'h02;
mem[16'h1A1D] = 8'h42;
mem[16'h1A1E] = 8'h3C;
mem[16'h1A1F] = 8'h00;
mem[16'h1A20] = 8'h3E;
mem[16'h1A21] = 8'h44;
mem[16'h1A22] = 8'h44;
mem[16'h1A23] = 8'h44;
mem[16'h1A24] = 8'h44;
mem[16'h1A25] = 8'h44;
mem[16'h1A26] = 8'h3E;
mem[16'h1A27] = 8'h00;
mem[16'h1A28] = 8'h7E;
mem[16'h1A29] = 8'h02;
mem[16'h1A2A] = 8'h02;
mem[16'h1A2B] = 8'h1E;
mem[16'h1A2C] = 8'h02;
mem[16'h1A2D] = 8'h02;
mem[16'h1A2E] = 8'h7E;
mem[16'h1A2F] = 8'h00;
mem[16'h1A30] = 8'h7E;
mem[16'h1A31] = 8'h02;
mem[16'h1A32] = 8'h02;
mem[16'h1A33] = 8'h1E;
mem[16'h1A34] = 8'h02;
mem[16'h1A35] = 8'h02;
mem[16'h1A36] = 8'h02;
mem[16'h1A37] = 8'h00;
mem[16'h1A38] = 8'h3C;
mem[16'h1A39] = 8'h42;
mem[16'h1A3A] = 8'h02;
mem[16'h1A3B] = 8'h72;
mem[16'h1A3C] = 8'h42;
mem[16'h1A3D] = 8'h42;
mem[16'h1A3E] = 8'h3C;
mem[16'h1A3F] = 8'h00;
mem[16'h1A40] = 8'h42;
mem[16'h1A41] = 8'h42;
mem[16'h1A42] = 8'h42;
mem[16'h1A43] = 8'h7E;
mem[16'h1A44] = 8'h42;
mem[16'h1A45] = 8'h42;
mem[16'h1A46] = 8'h42;
mem[16'h1A47] = 8'h00;
mem[16'h1A48] = 8'h38;
mem[16'h1A49] = 8'h10;
mem[16'h1A4A] = 8'h10;
mem[16'h1A4B] = 8'h10;
mem[16'h1A4C] = 8'h10;
mem[16'h1A4D] = 8'h10;
mem[16'h1A4E] = 8'h38;
mem[16'h1A4F] = 8'h00;
mem[16'h1A50] = 8'h70;
mem[16'h1A51] = 8'h20;
mem[16'h1A52] = 8'h20;
mem[16'h1A53] = 8'h20;
mem[16'h1A54] = 8'h20;
mem[16'h1A55] = 8'h22;
mem[16'h1A56] = 8'h1C;
mem[16'h1A57] = 8'h00;
mem[16'h1A58] = 8'h42;
mem[16'h1A59] = 8'h22;
mem[16'h1A5A] = 8'h12;
mem[16'h1A5B] = 8'h0E;
mem[16'h1A5C] = 8'h12;
mem[16'h1A5D] = 8'h22;
mem[16'h1A5E] = 8'h42;
mem[16'h1A5F] = 8'h00;
mem[16'h1A60] = 8'h02;
mem[16'h1A61] = 8'h02;
mem[16'h1A62] = 8'h02;
mem[16'h1A63] = 8'h02;
mem[16'h1A64] = 8'h02;
mem[16'h1A65] = 8'h02;
mem[16'h1A66] = 8'h7E;
mem[16'h1A67] = 8'h00;
mem[16'h1A68] = 8'h42;
mem[16'h1A69] = 8'h66;
mem[16'h1A6A] = 8'h5A;
mem[16'h1A6B] = 8'h5A;
mem[16'h1A6C] = 8'h42;
mem[16'h1A6D] = 8'h42;
mem[16'h1A6E] = 8'h42;
mem[16'h1A6F] = 8'h00;
mem[16'h1A70] = 8'h42;
mem[16'h1A71] = 8'h46;
mem[16'h1A72] = 8'h4A;
mem[16'h1A73] = 8'h52;
mem[16'h1A74] = 8'h62;
mem[16'h1A75] = 8'h42;
mem[16'h1A76] = 8'h42;
mem[16'h1A77] = 8'h00;
mem[16'h1A78] = 8'h3C;
mem[16'h1A79] = 8'h42;
mem[16'h1A7A] = 8'h42;
mem[16'h1A7B] = 8'h42;
mem[16'h1A7C] = 8'h42;
mem[16'h1A7D] = 8'h42;
mem[16'h1A7E] = 8'h3C;
mem[16'h1A7F] = 8'h00;
mem[16'h1A80] = 8'h3E;
mem[16'h1A81] = 8'h42;
mem[16'h1A82] = 8'h42;
mem[16'h1A83] = 8'h3E;
mem[16'h1A84] = 8'h02;
mem[16'h1A85] = 8'h02;
mem[16'h1A86] = 8'h02;
mem[16'h1A87] = 8'h00;
mem[16'h1A88] = 8'h3C;
mem[16'h1A89] = 8'h42;
mem[16'h1A8A] = 8'h42;
mem[16'h1A8B] = 8'h42;
mem[16'h1A8C] = 8'h52;
mem[16'h1A8D] = 8'h22;
mem[16'h1A8E] = 8'h5C;
mem[16'h1A8F] = 8'h00;
mem[16'h1A90] = 8'h3E;
mem[16'h1A91] = 8'h42;
mem[16'h1A92] = 8'h42;
mem[16'h1A93] = 8'h3E;
mem[16'h1A94] = 8'h12;
mem[16'h1A95] = 8'h22;
mem[16'h1A96] = 8'h42;
mem[16'h1A97] = 8'h00;
mem[16'h1A98] = 8'h3C;
mem[16'h1A99] = 8'h42;
mem[16'h1A9A] = 8'h02;
mem[16'h1A9B] = 8'h3C;
mem[16'h1A9C] = 8'h40;
mem[16'h1A9D] = 8'h42;
mem[16'h1A9E] = 8'h3C;
mem[16'h1A9F] = 8'h00;
mem[16'h1AA0] = 8'h7C;
mem[16'h1AA1] = 8'h10;
mem[16'h1AA2] = 8'h10;
mem[16'h1AA3] = 8'h10;
mem[16'h1AA4] = 8'h10;
mem[16'h1AA5] = 8'h10;
mem[16'h1AA6] = 8'h10;
mem[16'h1AA7] = 8'h00;
mem[16'h1AA8] = 8'h42;
mem[16'h1AA9] = 8'h42;
mem[16'h1AAA] = 8'h42;
mem[16'h1AAB] = 8'h42;
mem[16'h1AAC] = 8'h42;
mem[16'h1AAD] = 8'h42;
mem[16'h1AAE] = 8'h3C;
mem[16'h1AAF] = 8'h00;
mem[16'h1AB0] = 8'h42;
mem[16'h1AB1] = 8'h42;
mem[16'h1AB2] = 8'h42;
mem[16'h1AB3] = 8'h24;
mem[16'h1AB4] = 8'h24;
mem[16'h1AB5] = 8'h18;
mem[16'h1AB6] = 8'h18;
mem[16'h1AB7] = 8'h00;
mem[16'h1AB8] = 8'h42;
mem[16'h1AB9] = 8'h42;
mem[16'h1ABA] = 8'h42;
mem[16'h1ABB] = 8'h5A;
mem[16'h1ABC] = 8'h5A;
mem[16'h1ABD] = 8'h66;
mem[16'h1ABE] = 8'h42;
mem[16'h1ABF] = 8'h00;
mem[16'h1AC0] = 8'h42;
mem[16'h1AC1] = 8'h42;
mem[16'h1AC2] = 8'h24;
mem[16'h1AC3] = 8'h18;
mem[16'h1AC4] = 8'h24;
mem[16'h1AC5] = 8'h42;
mem[16'h1AC6] = 8'h42;
mem[16'h1AC7] = 8'h00;
mem[16'h1AC8] = 8'h44;
mem[16'h1AC9] = 8'h44;
mem[16'h1ACA] = 8'h44;
mem[16'h1ACB] = 8'h38;
mem[16'h1ACC] = 8'h10;
mem[16'h1ACD] = 8'h10;
mem[16'h1ACE] = 8'h10;
mem[16'h1ACF] = 8'h00;
mem[16'h1AD0] = 8'h7E;
mem[16'h1AD1] = 8'h40;
mem[16'h1AD2] = 8'h20;
mem[16'h1AD3] = 8'h18;
mem[16'h1AD4] = 8'h04;
mem[16'h1AD5] = 8'h02;
mem[16'h1AD6] = 8'h7E;
mem[16'h1AD7] = 8'h00;
mem[16'h1AD8] = 8'h3C;
mem[16'h1AD9] = 8'h04;
mem[16'h1ADA] = 8'h04;
mem[16'h1ADB] = 8'h04;
mem[16'h1ADC] = 8'h04;
mem[16'h1ADD] = 8'h04;
mem[16'h1ADE] = 8'h3C;
mem[16'h1ADF] = 8'h00;
mem[16'h1AE0] = 8'h00;
mem[16'h1AE1] = 8'h02;
mem[16'h1AE2] = 8'h04;
mem[16'h1AE3] = 8'h08;
mem[16'h1AE4] = 8'h10;
mem[16'h1AE5] = 8'h20;
mem[16'h1AE6] = 8'h40;
mem[16'h1AE7] = 8'h00;
mem[16'h1AE8] = 8'h3C;
mem[16'h1AE9] = 8'h20;
mem[16'h1AEA] = 8'h20;
mem[16'h1AEB] = 8'h20;
mem[16'h1AEC] = 8'h20;
mem[16'h1AED] = 8'h20;
mem[16'h1AEE] = 8'h3C;
mem[16'h1AEF] = 8'h00;
mem[16'h1AF0] = 8'h10;
mem[16'h1AF1] = 8'h28;
mem[16'h1AF2] = 8'h44;
mem[16'h1AF3] = 8'h00;
mem[16'h1AF4] = 8'h00;
mem[16'h1AF5] = 8'h00;
mem[16'h1AF6] = 8'h00;
mem[16'h1AF7] = 8'h00;
mem[16'h1AF8] = 8'h02;
mem[16'h1AF9] = 8'h00;
mem[16'h1AFA] = 8'h00;
mem[16'h1AFB] = 8'h00;
mem[16'h1AFC] = 8'h00;
mem[16'h1AFD] = 8'h00;
mem[16'h1AFE] = 8'h00;
mem[16'h1AFF] = 8'hFF;
mem[16'h1B00] = 8'h08;
mem[16'h1B01] = 8'h10;
mem[16'h1B02] = 8'h20;
mem[16'h1B03] = 8'h00;
mem[16'h1B04] = 8'h00;
mem[16'h1B05] = 8'h00;
mem[16'h1B06] = 8'h00;
mem[16'h1B07] = 8'h00;
mem[16'h1B08] = 8'h00;
mem[16'h1B09] = 8'h00;
mem[16'h1B0A] = 8'h1C;
mem[16'h1B0B] = 8'h20;
mem[16'h1B0C] = 8'h3C;
mem[16'h1B0D] = 8'h22;
mem[16'h1B0E] = 8'h5C;
mem[16'h1B0F] = 8'h00;
mem[16'h1B10] = 8'h02;
mem[16'h1B11] = 8'h02;
mem[16'h1B12] = 8'h3A;
mem[16'h1B13] = 8'h46;
mem[16'h1B14] = 8'h42;
mem[16'h1B15] = 8'h46;
mem[16'h1B16] = 8'h3A;
mem[16'h1B17] = 8'h00;
mem[16'h1B18] = 8'h00;
mem[16'h1B19] = 8'h00;
mem[16'h1B1A] = 8'h3C;
mem[16'h1B1B] = 8'h02;
mem[16'h1B1C] = 8'h02;
mem[16'h1B1D] = 8'h02;
mem[16'h1B1E] = 8'h3C;
mem[16'h1B1F] = 8'h00;
mem[16'h1B20] = 8'h40;
mem[16'h1B21] = 8'h40;
mem[16'h1B22] = 8'h5C;
mem[16'h1B23] = 8'h62;
mem[16'h1B24] = 8'h42;
mem[16'h1B25] = 8'h62;
mem[16'h1B26] = 8'h5C;
mem[16'h1B27] = 8'h00;
mem[16'h1B28] = 8'h00;
mem[16'h1B29] = 8'h00;
mem[16'h1B2A] = 8'h3C;
mem[16'h1B2B] = 8'h42;
mem[16'h1B2C] = 8'h7E;
mem[16'h1B2D] = 8'h02;
mem[16'h1B2E] = 8'h3C;
mem[16'h1B2F] = 8'h00;
mem[16'h1B30] = 8'h30;
mem[16'h1B31] = 8'h48;
mem[16'h1B32] = 8'h08;
mem[16'h1B33] = 8'h3E;
mem[16'h1B34] = 8'h08;
mem[16'h1B35] = 8'h08;
mem[16'h1B36] = 8'h08;
mem[16'h1B37] = 8'h00;
mem[16'h1B38] = 8'h00;
mem[16'h1B39] = 8'h00;
mem[16'h1B3A] = 8'h5C;
mem[16'h1B3B] = 8'h62;
mem[16'h1B3C] = 8'h62;
mem[16'h1B3D] = 8'h5C;
mem[16'h1B3E] = 8'h40;
mem[16'h1B3F] = 8'h3C;
mem[16'h1B40] = 8'h02;
mem[16'h1B41] = 8'h02;
mem[16'h1B42] = 8'h3A;
mem[16'h1B43] = 8'h46;
mem[16'h1B44] = 8'h42;
mem[16'h1B45] = 8'h42;
mem[16'h1B46] = 8'h42;
mem[16'h1B47] = 8'h00;
mem[16'h1B48] = 8'h10;
mem[16'h1B49] = 8'h00;
mem[16'h1B4A] = 8'h18;
mem[16'h1B4B] = 8'h10;
mem[16'h1B4C] = 8'h10;
mem[16'h1B4D] = 8'h10;
mem[16'h1B4E] = 8'h38;
mem[16'h1B4F] = 8'h00;
mem[16'h1B50] = 8'h20;
mem[16'h1B51] = 8'h00;
mem[16'h1B52] = 8'h30;
mem[16'h1B53] = 8'h20;
mem[16'h1B54] = 8'h20;
mem[16'h1B55] = 8'h20;
mem[16'h1B56] = 8'h22;
mem[16'h1B57] = 8'h1C;
mem[16'h1B58] = 8'h02;
mem[16'h1B59] = 8'h02;
mem[16'h1B5A] = 8'h22;
mem[16'h1B5B] = 8'h12;
mem[16'h1B5C] = 8'h0A;
mem[16'h1B5D] = 8'h16;
mem[16'h1B5E] = 8'h22;
mem[16'h1B5F] = 8'h00;
mem[16'h1B60] = 8'h18;
mem[16'h1B61] = 8'h10;
mem[16'h1B62] = 8'h10;
mem[16'h1B63] = 8'h10;
mem[16'h1B64] = 8'h10;
mem[16'h1B65] = 8'h10;
mem[16'h1B66] = 8'h38;
mem[16'h1B67] = 8'h00;
mem[16'h1B68] = 8'h00;
mem[16'h1B69] = 8'h00;
mem[16'h1B6A] = 8'h2E;
mem[16'h1B6B] = 8'h54;
mem[16'h1B6C] = 8'h54;
mem[16'h1B6D] = 8'h54;
mem[16'h1B6E] = 8'h54;
mem[16'h1B6F] = 8'h00;
mem[16'h1B70] = 8'h00;
mem[16'h1B71] = 8'h00;
mem[16'h1B72] = 8'h3E;
mem[16'h1B73] = 8'h44;
mem[16'h1B74] = 8'h44;
mem[16'h1B75] = 8'h44;
mem[16'h1B76] = 8'h44;
mem[16'h1B77] = 8'h00;
mem[16'h1B78] = 8'h00;
mem[16'h1B79] = 8'h00;
mem[16'h1B7A] = 8'h38;
mem[16'h1B7B] = 8'h44;
mem[16'h1B7C] = 8'h44;
mem[16'h1B7D] = 8'h44;
mem[16'h1B7E] = 8'h38;
mem[16'h1B7F] = 8'h00;
mem[16'h1B80] = 8'h00;
mem[16'h1B81] = 8'h00;
mem[16'h1B82] = 8'h3A;
mem[16'h1B83] = 8'h46;
mem[16'h1B84] = 8'h46;
mem[16'h1B85] = 8'h3A;
mem[16'h1B86] = 8'h02;
mem[16'h1B87] = 8'h02;
mem[16'h1B88] = 8'h00;
mem[16'h1B89] = 8'h00;
mem[16'h1B8A] = 8'h5C;
mem[16'h1B8B] = 8'h62;
mem[16'h1B8C] = 8'h62;
mem[16'h1B8D] = 8'h5C;
mem[16'h1B8E] = 8'h40;
mem[16'h1B8F] = 8'h40;
mem[16'h1B90] = 8'h00;
mem[16'h1B91] = 8'h00;
mem[16'h1B92] = 8'h3A;
mem[16'h1B93] = 8'h46;
mem[16'h1B94] = 8'h02;
mem[16'h1B95] = 8'h02;
mem[16'h1B96] = 8'h02;
mem[16'h1B97] = 8'h00;
mem[16'h1B98] = 8'h00;
mem[16'h1B99] = 8'h00;
mem[16'h1B9A] = 8'h7C;
mem[16'h1B9B] = 8'h02;
mem[16'h1B9C] = 8'h3C;
mem[16'h1B9D] = 8'h40;
mem[16'h1B9E] = 8'h3E;
mem[16'h1B9F] = 8'h00;
mem[16'h1BA0] = 8'h08;
mem[16'h1BA1] = 8'h08;
mem[16'h1BA2] = 8'h3E;
mem[16'h1BA3] = 8'h08;
mem[16'h1BA4] = 8'h08;
mem[16'h1BA5] = 8'h48;
mem[16'h1BA6] = 8'h30;
mem[16'h1BA7] = 8'h00;
mem[16'h1BA8] = 8'h00;
mem[16'h1BA9] = 8'h00;
mem[16'h1BAA] = 8'h42;
mem[16'h1BAB] = 8'h42;
mem[16'h1BAC] = 8'h42;
mem[16'h1BAD] = 8'h62;
mem[16'h1BAE] = 8'h5C;
mem[16'h1BAF] = 8'h00;
mem[16'h1BB0] = 8'h00;
mem[16'h1BB1] = 8'h00;
mem[16'h1BB2] = 8'h42;
mem[16'h1BB3] = 8'h42;
mem[16'h1BB4] = 8'h42;
mem[16'h1BB5] = 8'h24;
mem[16'h1BB6] = 8'h18;
mem[16'h1BB7] = 8'h00;
mem[16'h1BB8] = 8'h00;
mem[16'h1BB9] = 8'h00;
mem[16'h1BBA] = 8'h44;
mem[16'h1BBB] = 8'h44;
mem[16'h1BBC] = 8'h54;
mem[16'h1BBD] = 8'h54;
mem[16'h1BBE] = 8'h6C;
mem[16'h1BBF] = 8'h00;
mem[16'h1BC0] = 8'h00;
mem[16'h1BC1] = 8'h00;
mem[16'h1BC2] = 8'h42;
mem[16'h1BC3] = 8'h24;
mem[16'h1BC4] = 8'h18;
mem[16'h1BC5] = 8'h24;
mem[16'h1BC6] = 8'h42;
mem[16'h1BC7] = 8'h00;
mem[16'h1BC8] = 8'h00;
mem[16'h1BC9] = 8'h00;
mem[16'h1BCA] = 8'h42;
mem[16'h1BCB] = 8'h42;
mem[16'h1BCC] = 8'h62;
mem[16'h1BCD] = 8'h5C;
mem[16'h1BCE] = 8'h40;
mem[16'h1BCF] = 8'h3C;
mem[16'h1BD0] = 8'h00;
mem[16'h1BD1] = 8'h00;
mem[16'h1BD2] = 8'h7E;
mem[16'h1BD3] = 8'h20;
mem[16'h1BD4] = 8'h18;
mem[16'h1BD5] = 8'h04;
mem[16'h1BD6] = 8'h7E;
mem[16'h1BD7] = 8'h00;
mem[16'h1BD8] = 8'h38;
mem[16'h1BD9] = 8'h04;
mem[16'h1BDA] = 8'h04;
mem[16'h1BDB] = 8'h06;
mem[16'h1BDC] = 8'h04;
mem[16'h1BDD] = 8'h04;
mem[16'h1BDE] = 8'h38;
mem[16'h1BDF] = 8'h00;
mem[16'h1BE0] = 8'h08;
mem[16'h1BE1] = 8'h08;
mem[16'h1BE2] = 8'h08;
mem[16'h1BE3] = 8'h08;
mem[16'h1BE4] = 8'h08;
mem[16'h1BE5] = 8'h08;
mem[16'h1BE6] = 8'h08;
mem[16'h1BE7] = 8'h08;
mem[16'h1BE8] = 8'h0E;
mem[16'h1BE9] = 8'h10;
mem[16'h1BEA] = 8'h10;
mem[16'h1BEB] = 8'h30;
mem[16'h1BEC] = 8'h10;
mem[16'h1BED] = 8'h10;
mem[16'h1BEE] = 8'h0E;
mem[16'h1BEF] = 8'h00;
mem[16'h1BF0] = 8'h28;
mem[16'h1BF1] = 8'h14;
mem[16'h1BF2] = 8'h00;
mem[16'h1BF3] = 8'h00;
mem[16'h1BF4] = 8'h00;
mem[16'h1BF5] = 8'h00;
mem[16'h1BF6] = 8'h00;
mem[16'h1BF7] = 8'h00;
mem[16'h1BF8] = 8'hFF;
mem[16'h1BF9] = 8'hFF;
mem[16'h1BFA] = 8'hFF;
mem[16'h1BFB] = 8'hFF;
mem[16'h1BFC] = 8'hFF;
mem[16'h1BFD] = 8'h0F;
mem[16'h1BFE] = 8'hAB;
mem[16'h1BFF] = 8'h81;
mem[16'h1C00] = 8'h4C;
mem[16'h1C01] = 8'h5F;
mem[16'h1C02] = 8'h9C;
mem[16'h1C03] = 8'hA9;
mem[16'h1C04] = 8'h00;
mem[16'h1C05] = 8'h8D;
mem[16'h1C06] = 8'h06;
mem[16'h1C07] = 8'hA0;
mem[16'h1C08] = 8'h8D;
mem[16'h1C09] = 8'h09;
mem[16'h1C0A] = 8'hA0;
mem[16'h1C0B] = 8'h8D;
mem[16'h1C0C] = 8'h0A;
mem[16'h1C0D] = 8'hA0;
mem[16'h1C0E] = 8'hA9;
mem[16'h1C0F] = 8'h05;
mem[16'h1C10] = 8'h8D;
mem[16'h1C11] = 8'h07;
mem[16'h1C12] = 8'hA0;
mem[16'h1C13] = 8'hAD;
mem[16'h1C14] = 8'h19;
mem[16'h1C15] = 8'hA0;
mem[16'h1C16] = 8'hC9;
mem[16'h1C17] = 8'h1F;
mem[16'h1C18] = 8'hD0;
mem[16'h1C19] = 8'h1A;
mem[16'h1C1A] = 8'h10;
mem[16'h1C1B] = 8'h01;
mem[16'h1C1C] = 8'h85;
mem[16'h1C1D] = 8'hCD;
mem[16'h1C1E] = 8'h10;
mem[16'h1C1F] = 8'hC0;
mem[16'h1C20] = 8'hCE;
mem[16'h1C21] = 8'hF3;
mem[16'h1C22] = 8'h03;
mem[16'h1C23] = 8'hD0;
mem[16'h1C24] = 8'hFB;
mem[16'h1C25] = 8'hAD;
mem[16'h1C26] = 8'h00;
mem[16'h1C27] = 8'hC0;
mem[16'h1C28] = 8'h30;
mem[16'h1C29] = 8'h0A;
mem[16'h1C2A] = 8'hCE;
mem[16'h1C2B] = 8'hF4;
mem[16'h1C2C] = 8'h03;
mem[16'h1C2D] = 8'hD0;
mem[16'h1C2E] = 8'hF1;
mem[16'h1C2F] = 8'hCE;
mem[16'h1C30] = 8'h19;
mem[16'h1C31] = 8'hA0;
mem[16'h1C32] = 8'hD0;
mem[16'h1C33] = 8'hEC;
mem[16'h1C34] = 8'hA9;
mem[16'h1C35] = 8'h1F;
mem[16'h1C36] = 8'h8D;
mem[16'h1C37] = 8'h19;
mem[16'h1C38] = 8'hA0;
mem[16'h1C39] = 8'h20;
mem[16'h1C3A] = 8'h00;
mem[16'h1C3B] = 8'h0D;
mem[16'h1C3C] = 8'hEA;
mem[16'h1C3D] = 8'hEA;
mem[16'h1C3E] = 8'hA9;
mem[16'h1C3F] = 8'hFF;
mem[16'h1C40] = 8'h85;
mem[16'h1C41] = 8'h3A;
mem[16'h1C42] = 8'hA9;
mem[16'h1C43] = 8'hBF;
mem[16'h1C44] = 8'h85;
mem[16'h1C45] = 8'h3B;
mem[16'h1C46] = 8'hA0;
mem[16'h1C47] = 8'h13;
mem[16'h1C48] = 8'hD1;
mem[16'h1C49] = 8'h3A;
mem[16'h1C4A] = 8'hA0;
mem[16'h1C4B] = 8'h07;
mem[16'h1C4C] = 8'hB1;
mem[16'h1C4D] = 8'h3A;
mem[16'h1C4E] = 8'hC9;
mem[16'h1C4F] = 8'hA0;
mem[16'h1C50] = 8'hD0;
mem[16'h1C51] = 8'h02;
mem[16'h1C52] = 8'h60;
mem[16'h1C53] = 8'hA9;
mem[16'h1C54] = 8'hC9;
mem[16'h1C55] = 8'hC4;
mem[16'h1C56] = 8'hF0;
mem[16'h1C57] = 8'hFA;
mem[16'h1C58] = 8'hC9;
mem[16'h1C59] = 8'hCA;
mem[16'h1C5A] = 8'hF0;
mem[16'h1C5B] = 8'hF6;
mem[16'h1C5C] = 8'h4C;
mem[16'h1C5D] = 8'h4A;
mem[16'h1C5E] = 8'h9C;
mem[16'h1C5F] = 8'hA0;
mem[16'h1C60] = 8'h00;
mem[16'h1C61] = 8'h84;
mem[16'h1C62] = 8'h00;
mem[16'h1C63] = 8'h84;
mem[16'h1C64] = 8'h02;
mem[16'h1C65] = 8'hA9;
mem[16'h1C66] = 8'h97;
mem[16'h1C67] = 8'h85;
mem[16'h1C68] = 8'h01;
mem[16'h1C69] = 8'hA9;
mem[16'h1C6A] = 8'h03;
mem[16'h1C6B] = 8'h85;
mem[16'h1C6C] = 8'h03;
mem[16'h1C6D] = 8'hA2;
mem[16'h1C6E] = 8'h05;
mem[16'h1C6F] = 8'hAD;
mem[16'h1C70] = 8'h55;
mem[16'h1C71] = 8'hC0;
mem[16'h1C72] = 8'hEA;
mem[16'h1C73] = 8'hEA;
mem[16'h1C74] = 8'hEA;
mem[16'h1C75] = 8'hEA;
mem[16'h1C76] = 8'hEA;
mem[16'h1C77] = 8'hEA;
mem[16'h1C78] = 8'hEA;
mem[16'h1C79] = 8'hEA;
mem[16'h1C7A] = 8'hEA;
mem[16'h1C7B] = 8'hB1;
mem[16'h1C7C] = 8'h00;
mem[16'h1C7D] = 8'h91;
mem[16'h1C7E] = 8'h02;
mem[16'h1C7F] = 8'hC8;
mem[16'h1C80] = 8'hD0;
mem[16'h1C81] = 8'hF9;
mem[16'h1C82] = 8'hE6;
mem[16'h1C83] = 8'h01;
mem[16'h1C84] = 8'hE6;
mem[16'h1C85] = 8'h03;
mem[16'h1C86] = 8'hCA;
mem[16'h1C87] = 8'hD0;
mem[16'h1C88] = 8'hF2;
mem[16'h1C89] = 8'h4C;
mem[16'h1C8A] = 8'h03;
mem[16'h1C8B] = 8'h40;
mem[16'h1C8C] = 8'h84;
mem[16'h1C8D] = 8'hC2;
mem[16'h1C8E] = 8'hCC;
mem[16'h1C8F] = 8'hCF;
mem[16'h1C90] = 8'hED;
mem[16'h1C91] = 8'hFD;
mem[16'h1C92] = 8'h20;
mem[16'h1C93] = 8'h3A;
mem[16'h1C94] = 8'hFF;
mem[16'h1C95] = 8'hA9;
mem[16'h1C96] = 8'hA1;
mem[16'h1C97] = 8'h85;
mem[16'h1C98] = 8'h33;
mem[16'h1C99] = 8'h20;
mem[16'h1C9A] = 8'h67;
mem[16'h1C9B] = 8'hFD;
mem[16'h1C9C] = 8'h20;
mem[16'h1C9D] = 8'hC7;
mem[16'h1C9E] = 8'hFF;
mem[16'h1C9F] = 8'hAD;
mem[16'h1CA0] = 8'h00;
mem[16'h1CA1] = 8'h02;
mem[16'h1CA2] = 8'hC9;
mem[16'h1CA3] = 8'hA0;
mem[16'h1CA4] = 8'hF0;
mem[16'h1CA5] = 8'h13;
mem[16'h1CA6] = 8'hC8;
mem[16'h1CA7] = 8'hC9;
mem[16'h1CA8] = 8'hA4;
mem[16'h1CA9] = 8'hF0;
mem[16'h1CAA] = 8'h92;
mem[16'h1CAB] = 8'h88;
mem[16'h1CAC] = 8'h20;
mem[16'h1CAD] = 8'hA7;
mem[16'h1CAE] = 8'hFF;
mem[16'h1CAF] = 8'hC9;
mem[16'h1CB0] = 8'h93;
mem[16'h1CB1] = 8'hD0;
mem[16'h1CB2] = 8'hD5;
mem[16'h1CB3] = 8'h8A;
mem[16'h1CB4] = 8'hF0;
mem[16'h1CB5] = 8'hD2;
mem[16'h1CB6] = 8'h20;
mem[16'h1CB7] = 8'h78;
mem[16'h1CB8] = 8'hFE;
mem[16'h1CB9] = 8'hA9;
mem[16'h1CBA] = 8'h03;
mem[16'h1CBB] = 8'h85;
mem[16'h1CBC] = 8'h3D;
mem[16'h1CBD] = 8'h20;
mem[16'h1CBE] = 8'h34;
mem[16'h1CBF] = 8'hF6;
mem[16'h1CC0] = 8'h0A;
mem[16'h1CC1] = 8'hE9;
mem[16'h1CC2] = 8'hBE;
mem[16'h1CC3] = 8'hC9;
mem[16'h1CC4] = 8'hC2;
mem[16'h1CC5] = 8'h90;
mem[16'h1CC6] = 8'hC1;
mem[16'h1CC7] = 8'h0A;
mem[16'h1CC8] = 8'h0A;
mem[16'h1CC9] = 8'hA2;
mem[16'h1CCA] = 8'h04;
mem[16'h1CCB] = 8'h0A;
mem[16'h1CCC] = 8'h26;
mem[16'h1CCD] = 8'h42;
mem[16'h1CCE] = 8'h26;
mem[16'h1CCF] = 8'h43;
mem[16'h1CD0] = 8'hCA;
mem[16'h1CD1] = 8'h10;
mem[16'h1CD2] = 8'hF8;
mem[16'h1CD3] = 8'hC6;
mem[16'h1CD4] = 8'h3D;
mem[16'h1CD5] = 8'hF0;
mem[16'h1CD6] = 8'hF4;
mem[16'h1CD7] = 8'h10;
mem[16'h1CD8] = 8'hE4;
mem[16'h1CD9] = 8'hA2;
mem[16'h1CDA] = 8'h05;
mem[16'h1CDB] = 8'h20;
mem[16'h1CDC] = 8'h34;
mem[16'h1CDD] = 8'hF6;
mem[16'h1CDE] = 8'h84;
mem[16'h1CDF] = 8'h34;
mem[16'h1CE0] = 8'hDD;
mem[16'h1CE1] = 8'hB4;
mem[16'h1CE2] = 8'hF9;
mem[16'h1CE3] = 8'hD0;
mem[16'h1CE4] = 8'h13;
mem[16'h1CE5] = 8'h20;
mem[16'h1CE6] = 8'h34;
mem[16'h1CE7] = 8'hF6;
mem[16'h1CE8] = 8'hDD;
mem[16'h1CE9] = 8'hBA;
mem[16'h1CEA] = 8'hF9;
mem[16'h1CEB] = 8'hF0;
mem[16'h1CEC] = 8'h0D;
mem[16'h1CED] = 8'hBD;
mem[16'h1CEE] = 8'hBA;
mem[16'h1CEF] = 8'hF9;
mem[16'h1CF0] = 8'hF0;
mem[16'h1CF1] = 8'h07;
mem[16'h1CF2] = 8'hC9;
mem[16'h1CF3] = 8'hA4;
mem[16'h1CF4] = 8'hF0;
mem[16'h1CF5] = 8'h03;
mem[16'h1CF6] = 8'hA4;
mem[16'h1CF7] = 8'h34;
mem[16'h1CF8] = 8'h18;
mem[16'h1CF9] = 8'h88;
mem[16'h1CFA] = 8'h26;
mem[16'h1CFB] = 8'h44;
mem[16'h1CFC] = 8'hE0;
mem[16'h1CFD] = 8'h03;
mem[16'h1CFE] = 8'hD0;
mem[16'h1CFF] = 8'h0D;
mem[16'h1D00] = 8'hB3;
mem[16'h1D01] = 8'hBD;
mem[16'h1D02] = 8'hC8;
mem[16'h1D03] = 8'hB4;
mem[16'h1D04] = 8'h29;
mem[16'h1D05] = 8'h7F;
mem[16'h1D06] = 8'h0D;
mem[16'h1D07] = 8'h9E;
mem[16'h1D08] = 8'hB3;
mem[16'h1D09] = 8'h9D;
mem[16'h1D0A] = 8'hC8;
mem[16'h1D0B] = 8'hB4;
mem[16'h1D0C] = 8'h20;
mem[16'h1D0D] = 8'h37;
mem[16'h1D0E] = 8'hB0;
mem[16'h1D0F] = 8'h4C;
mem[16'h1D10] = 8'h7F;
mem[16'h1D11] = 8'hB3;
mem[16'h1D12] = 8'h20;
mem[16'h1D13] = 8'h00;
mem[16'h1D14] = 8'hB3;
mem[16'h1D15] = 8'h4C;
mem[16'h1D16] = 8'h7F;
mem[16'h1D17] = 8'hB3;
mem[16'h1D18] = 8'h20;
mem[16'h1D19] = 8'h28;
mem[16'h1D1A] = 8'hAB;
mem[16'h1D1B] = 8'h20;
mem[16'h1D1C] = 8'hB6;
mem[16'h1D1D] = 8'hB0;
mem[16'h1D1E] = 8'hB0;
mem[16'h1D1F] = 8'hEF;
mem[16'h1D20] = 8'hEE;
mem[16'h1D21] = 8'hE4;
mem[16'h1D22] = 8'hB5;
mem[16'h1D23] = 8'hD0;
mem[16'h1D24] = 8'hF6;
mem[16'h1D25] = 8'hEE;
mem[16'h1D26] = 8'hE5;
mem[16'h1D27] = 8'hB5;
mem[16'h1D28] = 8'h4C;
mem[16'h1D29] = 8'h1B;
mem[16'h1D2A] = 8'hAD;
mem[16'h1D2B] = 8'h20;
mem[16'h1D2C] = 8'h28;
mem[16'h1D2D] = 8'hAB;
mem[16'h1D2E] = 8'hAE;
mem[16'h1D2F] = 8'h9C;
mem[16'h1D30] = 8'hB3;
mem[16'h1D31] = 8'hBD;
mem[16'h1D32] = 8'hC8;
mem[16'h1D33] = 8'hB4;
mem[16'h1D34] = 8'h10;
mem[16'h1D35] = 8'h03;
mem[16'h1D36] = 8'h4C;
mem[16'h1D37] = 8'h7B;
mem[16'h1D38] = 8'hB3;
mem[16'h1D39] = 8'hAE;
mem[16'h1D3A] = 8'h9C;
mem[16'h1D3B] = 8'hB3;
mem[16'h1D3C] = 8'hBD;
mem[16'h1D3D] = 8'hC6;
mem[16'h1D3E] = 8'hB4;
mem[16'h1D3F] = 8'h8D;
mem[16'h1D40] = 8'hD1;
mem[16'h1D41] = 8'hB5;
mem[16'h1D42] = 8'h9D;
mem[16'h1D43] = 8'hE6;
mem[16'h1D44] = 8'hB4;
mem[16'h1D45] = 8'hA9;
mem[16'h1D46] = 8'hFF;
mem[16'h1D47] = 8'h9D;
mem[16'h1D48] = 8'hC6;
mem[16'h1D49] = 8'hB4;
mem[16'h1D4A] = 8'hBC;
mem[16'h1D4B] = 8'hC7;
mem[16'h1D4C] = 8'hB4;
mem[16'h1D4D] = 8'h8C;
mem[16'h1D4E] = 8'hD2;
mem[16'h1D4F] = 8'hB5;
mem[16'h1D50] = 8'h20;
mem[16'h1D51] = 8'h37;
mem[16'h1D52] = 8'hB0;
mem[16'h1D53] = 8'h18;
mem[16'h1D54] = 8'h20;
mem[16'h1D55] = 8'h5E;
mem[16'h1D56] = 8'hAF;
mem[16'h1D57] = 8'hB0;
mem[16'h1D58] = 8'h2A;
mem[16'h1D59] = 8'h20;
mem[16'h1D5A] = 8'h0C;
mem[16'h1D5B] = 8'hAF;
mem[16'h1D5C] = 8'hA0;
mem[16'h1D5D] = 8'h0C;
mem[16'h1D5E] = 8'h8C;
mem[16'h1D5F] = 8'h9C;
mem[16'h1D60] = 8'hB3;
mem[16'h1D61] = 8'hB1;
mem[16'h1D62] = 8'h42;
mem[16'h1D63] = 8'h30;
mem[16'h1D64] = 8'h0B;
mem[16'h1D65] = 8'hF0;
mem[16'h1D66] = 8'h09;
mem[16'h1D67] = 8'h48;
mem[16'h1D68] = 8'hC8;
mem[16'h1D69] = 8'hB1;
mem[16'h1D6A] = 8'h42;
mem[16'h1D6B] = 8'hA8;
mem[16'h1D6C] = 8'h68;
mem[16'h1D6D] = 8'h20;
mem[16'h1D6E] = 8'h89;
mem[16'h1D6F] = 8'hAD;
mem[16'h1D70] = 8'hAC;
mem[16'h1D71] = 8'h9C;
mem[16'h1D72] = 8'hB3;
mem[16'h1D73] = 8'hC8;
mem[16'h1D74] = 8'hC8;
mem[16'h1D75] = 8'hD0;
mem[16'h1D76] = 8'hE7;
mem[16'h1D77] = 8'hAD;
mem[16'h1D78] = 8'hD3;
mem[16'h1D79] = 8'hB5;
mem[16'h1D7A] = 8'hAC;
mem[16'h1D7B] = 8'hD4;
mem[16'h1D7C] = 8'hB5;
mem[16'h1D7D] = 8'h20;
mem[16'h1D7E] = 8'h89;
mem[16'h1D7F] = 8'hAD;
mem[16'h1D80] = 8'h38;
mem[16'h1D81] = 8'hB0;
mem[16'h1D82] = 8'hD1;
mem[16'h1D83] = 8'h20;
mem[16'h1D84] = 8'hFB;
mem[16'h1D85] = 8'hAF;
mem[16'h1D86] = 8'h4C;
mem[16'h1D87] = 8'h7F;
mem[16'h1D88] = 8'hB3;
mem[16'h1D89] = 8'h38;
mem[16'h1D8A] = 8'h20;
mem[16'h1D8B] = 8'hDD;
mem[16'h1D8C] = 8'hB2;
mem[16'h1D8D] = 8'hA9;
mem[16'h1D8E] = 8'h00;
mem[16'h1D8F] = 8'hA2;
mem[16'h1D90] = 8'h05;
mem[16'h1D91] = 8'h9D;
mem[16'h1D92] = 8'hF0;
mem[16'h1D93] = 8'hB5;
mem[16'h1D94] = 8'hCA;
mem[16'h1D95] = 8'h10;
mem[16'h1D96] = 8'hFA;
mem[16'h1D97] = 8'h60;
mem[16'h1D98] = 8'h20;
mem[16'h1D99] = 8'hDC;
mem[16'h1D9A] = 8'hAB;
mem[16'h1D9B] = 8'hA9;
mem[16'h1D9C] = 8'hFF;
mem[16'h1D9D] = 8'h8D;
mem[16'h1D9E] = 8'hF9;
mem[16'h1D9F] = 8'hB5;
mem[16'h1DA0] = 8'h20;
mem[16'h1DA1] = 8'hF7;
mem[16'h1DA2] = 8'hAF;
mem[16'h1DA3] = 8'hA9;
mem[16'h1DA4] = 8'h16;
mem[16'h1DA5] = 8'h8D;
mem[16'h1DA6] = 8'h9D;
mem[16'h1DA7] = 8'hB3;
mem[16'h1DA8] = 8'h20;
mem[16'h1DA9] = 8'h2F;
mem[16'h1DAA] = 8'hAE;
mem[16'h1DAB] = 8'h20;
mem[16'h1DAC] = 8'h2F;
mem[16'h1DAD] = 8'hAE;
mem[16'h1DAE] = 8'hA2;
mem[16'h1DAF] = 8'h0B;
mem[16'h1DB0] = 8'hBD;
mem[16'h1DB1] = 8'hAF;
mem[16'h1DB2] = 8'hB3;
mem[16'h1DB3] = 8'h20;
mem[16'h1DB4] = 8'hED;
mem[16'h1DB5] = 8'hFD;
mem[16'h1DB6] = 8'hCA;
mem[16'h1DB7] = 8'h10;
mem[16'h1DB8] = 8'hF7;
mem[16'h1DB9] = 8'h86;
mem[16'h1DBA] = 8'h45;
mem[16'h1DBB] = 8'hAD;
mem[16'h1DBC] = 8'hF6;
mem[16'h1DBD] = 8'hB7;
mem[16'h1DBE] = 8'h85;
mem[16'h1DBF] = 8'h44;
mem[16'h1DC0] = 8'h20;
mem[16'h1DC1] = 8'h42;
mem[16'h1DC2] = 8'hAE;
mem[16'h1DC3] = 8'h20;
mem[16'h1DC4] = 8'h2F;
mem[16'h1DC5] = 8'hAE;
mem[16'h1DC6] = 8'h20;
mem[16'h1DC7] = 8'h2F;
mem[16'h1DC8] = 8'hAE;
mem[16'h1DC9] = 8'h18;
mem[16'h1DCA] = 8'h20;
mem[16'h1DCB] = 8'h11;
mem[16'h1DCC] = 8'hB0;
mem[16'h1DCD] = 8'hB0;
mem[16'h1DCE] = 8'h5D;
mem[16'h1DCF] = 8'hA2;
mem[16'h1DD0] = 8'h00;
mem[16'h1DD1] = 8'h8E;
mem[16'h1DD2] = 8'h9C;
mem[16'h1DD3] = 8'hB3;
mem[16'h1DD4] = 8'hBD;
mem[16'h1DD5] = 8'hC6;
mem[16'h1DD6] = 8'hB4;
mem[16'h1DD7] = 8'hF0;
mem[16'h1DD8] = 8'h53;
mem[16'h1DD9] = 8'h30;
mem[16'h1DDA] = 8'h4A;
mem[16'h1DDB] = 8'hA0;
mem[16'h1DDC] = 8'hA0;
mem[16'h1DDD] = 8'hBD;
mem[16'h1DDE] = 8'hC8;
mem[16'h1DDF] = 8'hB4;
mem[16'h1DE0] = 8'h10;
mem[16'h1DE1] = 8'h02;
mem[16'h1DE2] = 8'hA0;
mem[16'h1DE3] = 8'hAA;
mem[16'h1DE4] = 8'h98;
mem[16'h1DE5] = 8'h20;
mem[16'h1DE6] = 8'hED;
mem[16'h1DE7] = 8'hFD;
mem[16'h1DE8] = 8'hBD;
mem[16'h1DE9] = 8'hC8;
mem[16'h1DEA] = 8'hB4;
mem[16'h1DEB] = 8'h29;
mem[16'h1DEC] = 8'h7F;
mem[16'h1DED] = 8'hA0;
mem[16'h1DEE] = 8'h07;
mem[16'h1DEF] = 8'h0A;
mem[16'h1DF0] = 8'h0A;
mem[16'h1DF1] = 8'hB0;
mem[16'h1DF2] = 8'h03;
mem[16'h1DF3] = 8'h88;
mem[16'h1DF4] = 8'hD0;
mem[16'h1DF5] = 8'hFA;
mem[16'h1DF6] = 8'hB9;
mem[16'h1DF7] = 8'hA7;
mem[16'h1DF8] = 8'hB3;
mem[16'h1DF9] = 8'h20;
mem[16'h1DFA] = 8'hED;
mem[16'h1DFB] = 8'hFD;
mem[16'h1DFC] = 8'hA9;
mem[16'h1DFD] = 8'hA0;
mem[16'h1DFE] = 8'h20;
mem[16'h1DFF] = 8'hED;
mem[16'h1E00] = 8'hFD;
mem[16'h1E01] = 8'hBD;
mem[16'h1E02] = 8'hE7;
mem[16'h1E03] = 8'hB4;
mem[16'h1E04] = 8'h85;
mem[16'h1E05] = 8'h44;
mem[16'h1E06] = 8'hBD;
mem[16'h1E07] = 8'hE8;
mem[16'h1E08] = 8'hB4;
mem[16'h1E09] = 8'h85;
mem[16'h1E0A] = 8'h45;
mem[16'h1E0B] = 8'h20;
mem[16'h1E0C] = 8'h42;
mem[16'h1E0D] = 8'hAE;
mem[16'h1E0E] = 8'hA9;
mem[16'h1E0F] = 8'hA0;
mem[16'h1E10] = 8'h20;
mem[16'h1E11] = 8'hED;
mem[16'h1E12] = 8'hFD;
mem[16'h1E13] = 8'hE8;
mem[16'h1E14] = 8'hE8;
mem[16'h1E15] = 8'hE8;
mem[16'h1E16] = 8'hA0;
mem[16'h1E17] = 8'h1D;
mem[16'h1E18] = 8'hBD;
mem[16'h1E19] = 8'hC6;
mem[16'h1E1A] = 8'hB4;
mem[16'h1E1B] = 8'h20;
mem[16'h1E1C] = 8'hED;
mem[16'h1E1D] = 8'hFD;
mem[16'h1E1E] = 8'hE8;
mem[16'h1E1F] = 8'h88;
mem[16'h1E20] = 8'h10;
mem[16'h1E21] = 8'hF6;
mem[16'h1E22] = 8'h20;
mem[16'h1E23] = 8'h2F;
mem[16'h1E24] = 8'hAE;
mem[16'h1E25] = 8'h20;
mem[16'h1E26] = 8'h30;
mem[16'h1E27] = 8'hB2;
mem[16'h1E28] = 8'h90;
mem[16'h1E29] = 8'hA7;
mem[16'h1E2A] = 8'hB0;
mem[16'h1E2B] = 8'h9E;
mem[16'h1E2C] = 8'h4C;
mem[16'h1E2D] = 8'h7F;
mem[16'h1E2E] = 8'hB3;
mem[16'h1E2F] = 8'hA9;
mem[16'h1E30] = 8'h8D;
mem[16'h1E31] = 8'h20;
mem[16'h1E32] = 8'hED;
mem[16'h1E33] = 8'hFD;
mem[16'h1E34] = 8'hCE;
mem[16'h1E35] = 8'h9D;
mem[16'h1E36] = 8'hB3;
mem[16'h1E37] = 8'hD0;
mem[16'h1E38] = 8'h08;
mem[16'h1E39] = 8'h20;
mem[16'h1E3A] = 8'h0C;
mem[16'h1E3B] = 8'hFD;
mem[16'h1E3C] = 8'hA9;
mem[16'h1E3D] = 8'h15;
mem[16'h1E3E] = 8'h8D;
mem[16'h1E3F] = 8'h9D;
mem[16'h1E40] = 8'hB3;
mem[16'h1E41] = 8'h60;
mem[16'h1E42] = 8'hA0;
mem[16'h1E43] = 8'h02;
mem[16'h1E44] = 8'hA9;
mem[16'h1E45] = 8'h00;
mem[16'h1E46] = 8'h48;
mem[16'h1E47] = 8'hA5;
mem[16'h1E48] = 8'h44;
mem[16'h1E49] = 8'hD9;
mem[16'h1E4A] = 8'hA4;
mem[16'h1E4B] = 8'hB3;
mem[16'h1E4C] = 8'h90;
mem[16'h1E4D] = 8'h12;
mem[16'h1E4E] = 8'hF9;
mem[16'h1E4F] = 8'hA4;
mem[16'h1E50] = 8'hB3;
mem[16'h1E51] = 8'h85;
mem[16'h1E52] = 8'h44;
mem[16'h1E53] = 8'hA5;
mem[16'h1E54] = 8'h45;
mem[16'h1E55] = 8'hE9;
mem[16'h1E56] = 8'h00;
mem[16'h1E57] = 8'h85;
mem[16'h1E58] = 8'h45;
mem[16'h1E59] = 8'h68;
mem[16'h1E5A] = 8'h69;
mem[16'h1E5B] = 8'h00;
mem[16'h1E5C] = 8'h48;
mem[16'h1E5D] = 8'h4C;
mem[16'h1E5E] = 8'h47;
mem[16'h1E5F] = 8'hAE;
mem[16'h1E60] = 8'h68;
mem[16'h1E61] = 8'h09;
mem[16'h1E62] = 8'hB0;
mem[16'h1E63] = 8'h20;
mem[16'h1E64] = 8'hED;
mem[16'h1E65] = 8'hFD;
mem[16'h1E66] = 8'h88;
mem[16'h1E67] = 8'h10;
mem[16'h1E68] = 8'hDB;
mem[16'h1E69] = 8'h60;
mem[16'h1E6A] = 8'h20;
mem[16'h1E6B] = 8'h08;
mem[16'h1E6C] = 8'hAF;
mem[16'h1E6D] = 8'hA0;
mem[16'h1E6E] = 8'h00;
mem[16'h1E6F] = 8'h8C;
mem[16'h1E70] = 8'hC5;
mem[16'h1E71] = 8'hB5;
mem[16'h1E72] = 8'hB1;
mem[16'h1E73] = 8'h42;
mem[16'h1E74] = 8'h99;
mem[16'h1E75] = 8'hD1;
mem[16'h1E76] = 8'hB5;
mem[16'h1E77] = 8'hC8;
mem[16'h1E78] = 8'hC0;
mem[16'h1E79] = 8'h2D;
mem[16'h1E7A] = 8'hD0;
mem[16'h1E7B] = 8'hF6;
mem[16'h1E7C] = 8'h18;
mem[16'h1E7D] = 8'h60;
mem[16'h1E7E] = 8'h20;
mem[16'h1E7F] = 8'h08;
mem[16'h1E80] = 8'hAF;
mem[16'h1E81] = 8'hA0;
mem[16'h1E82] = 8'h00;
mem[16'h1E83] = 8'hB9;
mem[16'h1E84] = 8'hD1;
mem[16'h1E85] = 8'hB5;
mem[16'h1E86] = 8'h91;
mem[16'h1E87] = 8'h42;
mem[16'h1E88] = 8'hC8;
mem[16'h1E89] = 8'hC0;
mem[16'h1E8A] = 8'h2D;
mem[16'h1E8B] = 8'hD0;
mem[16'h1E8C] = 8'hF6;
mem[16'h1E8D] = 8'h60;
mem[16'h1E8E] = 8'h20;
mem[16'h1E8F] = 8'hDC;
mem[16'h1E90] = 8'hAB;
mem[16'h1E91] = 8'hA9;
mem[16'h1E92] = 8'h04;
mem[16'h1E93] = 8'h20;
mem[16'h1E94] = 8'h58;
mem[16'h1E95] = 8'hB0;
mem[16'h1E96] = 8'hAD;
mem[16'h1E97] = 8'hF9;
mem[16'h1E98] = 8'hB5;
mem[16'h1E99] = 8'h49;
mem[16'h1E9A] = 8'hFF;
mem[16'h1E9B] = 8'h8D;
mem[16'h1E9C] = 8'hC1;
mem[16'h1E9D] = 8'hB3;
mem[16'h1E9E] = 8'hA9;
mem[16'h1E9F] = 8'h11;
mem[16'h1EA0] = 8'h8D;
mem[16'h1EA1] = 8'hEB;
mem[16'h1EA2] = 8'hB3;
mem[16'h1EA3] = 8'hA9;
mem[16'h1EA4] = 8'h01;
mem[16'h1EA5] = 8'h8D;
mem[16'h1EA6] = 8'hEC;
mem[16'h1EA7] = 8'hB3;
mem[16'h1EA8] = 8'hA2;
mem[16'h1EA9] = 8'h38;
mem[16'h1EAA] = 8'hA9;
mem[16'h1EAB] = 8'h00;
mem[16'h1EAC] = 8'h9D;
mem[16'h1EAD] = 8'hBB;
mem[16'h1EAE] = 8'hB3;
mem[16'h1EAF] = 8'hE8;
mem[16'h1EB0] = 8'hD0;
mem[16'h1EB1] = 8'hFA;
mem[16'h1EB2] = 8'hA2;
mem[16'h1EB3] = 8'h0C;
mem[16'h1EB4] = 8'hE0;
mem[16'h1EB5] = 8'h8C;
mem[16'h1EB6] = 8'hF0;
mem[16'h1EB7] = 8'h14;
mem[16'h1EB8] = 8'hA0;
mem[16'h1EB9] = 8'h03;
mem[16'h1EBA] = 8'hB9;
mem[16'h1EBB] = 8'hA0;
mem[16'h1EBC] = 8'hB3;
mem[16'h1EBD] = 8'h9D;
mem[16'h1EBE] = 8'hF3;
mem[16'h1EBF] = 8'hB3;
mem[16'h1EC0] = 8'hE8;
mem[16'h1EC1] = 8'h88;
mem[16'h1EC2] = 8'h10;
mem[16'h1EC3] = 8'hF6;
mem[16'h1EC4] = 8'hE0;
mem[16'h1EC5] = 8'h44;
mem[16'h1EC6] = 8'hD0;
mem[16'h1EC7] = 8'hEC;
mem[16'h1EC8] = 8'hA2;
mem[16'h1EC9] = 8'h48;
mem[16'h1ECA] = 8'hD0;
mem[16'h1ECB] = 8'hE8;
mem[16'h1ECC] = 8'h20;
mem[16'h1ECD] = 8'hFB;
mem[16'h1ECE] = 8'hAF;
mem[16'h1ECF] = 8'hA2;
mem[16'h1ED0] = 8'h00;
mem[16'h1ED1] = 8'h8A;
mem[16'h1ED2] = 8'h9D;
mem[16'h1ED3] = 8'hBB;
mem[16'h1ED4] = 8'hB4;
mem[16'h1ED5] = 8'hE8;
mem[16'h1ED6] = 8'hD0;
mem[16'h1ED7] = 8'hFA;
mem[16'h1ED8] = 8'h20;
mem[16'h1ED9] = 8'h45;
mem[16'h1EDA] = 8'hB0;
mem[16'h1EDB] = 8'hA9;
mem[16'h1EDC] = 8'h11;
mem[16'h1EDD] = 8'hAC;
mem[16'h1EDE] = 8'hF0;
mem[16'h1EDF] = 8'hB3;
mem[16'h1EE0] = 8'h88;
mem[16'h1EE1] = 8'h88;
mem[16'h1EE2] = 8'h8D;
mem[16'h1EE3] = 8'hEC;
mem[16'h1EE4] = 8'hB7;
mem[16'h1EE5] = 8'h8D;
mem[16'h1EE6] = 8'hBC;
mem[16'h1EE7] = 8'hB4;
mem[16'h1EE8] = 8'h8C;
mem[16'h1EE9] = 8'hBD;
mem[16'h1EEA] = 8'hB4;
mem[16'h1EEB] = 8'hC8;
mem[16'h1EEC] = 8'h8C;
mem[16'h1EED] = 8'hED;
mem[16'h1EEE] = 8'hB7;
mem[16'h1EEF] = 8'hA9;
mem[16'h1EF0] = 8'h02;
mem[16'h1EF1] = 8'h20;
mem[16'h1EF2] = 8'h58;
mem[16'h1EF3] = 8'hB0;
mem[16'h1EF4] = 8'hAC;
mem[16'h1EF5] = 8'hBD;
mem[16'h1EF6] = 8'hB4;
mem[16'h1EF7] = 8'h88;
mem[16'h1EF8] = 8'h30;
mem[16'h1EF9] = 8'h05;
mem[16'h1EFA] = 8'hD0;
mem[16'h1EFB] = 8'hEC;
mem[16'h1EFC] = 8'h98;
mem[16'h1EFD] = 8'hF0;
mem[16'h1EFE] = 8'hE6;
mem[16'h1EFF] = 8'h20;
mem[16'h1F00] = 8'hC2;
mem[16'h1F01] = 8'hB7;
mem[16'h1F02] = 8'h20;
mem[16'h1F03] = 8'h4A;
mem[16'h1F04] = 8'hB7;
mem[16'h1F05] = 8'h4C;
mem[16'h1F06] = 8'h7F;
mem[16'h1F07] = 8'hB3;
mem[16'h1F08] = 8'hA2;
mem[16'h1F09] = 8'h00;
mem[16'h1F0A] = 8'hF0;
mem[16'h1F0B] = 8'h06;
mem[16'h1F0C] = 8'hA2;
mem[16'h1F0D] = 8'h02;
mem[16'h1F0E] = 8'hD0;
mem[16'h1F0F] = 8'h02;
mem[16'h1F10] = 8'hA2;
mem[16'h1F11] = 8'h04;
mem[16'h1F12] = 8'hBD;
mem[16'h1F13] = 8'hC7;
mem[16'h1F14] = 8'hB5;
mem[16'h1F15] = 8'h85;
mem[16'h1F16] = 8'h42;
mem[16'h1F17] = 8'hBD;
mem[16'h1F18] = 8'hC8;
mem[16'h1F19] = 8'hB5;
mem[16'h1F1A] = 8'h85;
mem[16'h1F1B] = 8'h43;
mem[16'h1F1C] = 8'h60;
mem[16'h1F1D] = 8'h2C;
mem[16'h1F1E] = 8'hD5;
mem[16'h1F1F] = 8'hB5;
mem[16'h1F20] = 8'h70;
mem[16'h1F21] = 8'h01;
mem[16'h1F22] = 8'h60;
mem[16'h1F23] = 8'h20;
mem[16'h1F24] = 8'hE4;
mem[16'h1F25] = 8'hAF;
mem[16'h1F26] = 8'hA9;
mem[16'h1F27] = 8'h02;
mem[16'h1F28] = 8'h20;
mem[16'h1F29] = 8'h52;
mem[16'h1F2A] = 8'hB0;
mem[16'h1F2B] = 8'hA9;
mem[16'h1F2C] = 8'hBF;
mem[16'h1F2D] = 8'h2D;
mem[16'h1F2E] = 8'hD5;
mem[16'h1F2F] = 8'hB5;
mem[16'h1F30] = 8'h8D;
mem[16'h1F31] = 8'hD5;
mem[16'h1F32] = 8'hB5;
mem[16'h1F33] = 8'h60;
mem[16'h1F34] = 8'hAD;
mem[16'h1F35] = 8'hD5;
mem[16'h1F36] = 8'hB5;
mem[16'h1F37] = 8'h30;
mem[16'h1F38] = 8'h01;
mem[16'h1F39] = 8'h60;
mem[16'h1F3A] = 8'h20;
mem[16'h1F3B] = 8'h4B;
mem[16'h1F3C] = 8'hAF;
mem[16'h1F3D] = 8'hA9;
mem[16'h1F3E] = 8'h02;
mem[16'h1F3F] = 8'h20;
mem[16'h1F40] = 8'h52;
mem[16'h1F41] = 8'hB0;
mem[16'h1F42] = 8'hA9;
mem[16'h1F43] = 8'h7F;
mem[16'h1F44] = 8'h2D;
mem[16'h1F45] = 8'hD5;
mem[16'h1F46] = 8'hB5;
mem[16'h1F47] = 8'h8D;
mem[16'h1F48] = 8'hD5;
mem[16'h1F49] = 8'hB5;
mem[16'h1F4A] = 8'h60;
mem[16'h1F4B] = 8'hAD;
mem[16'h1F4C] = 8'hC9;
mem[16'h1F4D] = 8'hB5;
mem[16'h1F4E] = 8'h8D;
mem[16'h1F4F] = 8'hF0;
mem[16'h1F50] = 8'hB7;
mem[16'h1F51] = 8'hAD;
mem[16'h1F52] = 8'hCA;
mem[16'h1F53] = 8'hB5;
mem[16'h1F54] = 8'h8D;
mem[16'h1F55] = 8'hF1;
mem[16'h1F56] = 8'hB7;
mem[16'h1F57] = 8'hAE;
mem[16'h1F58] = 8'hD3;
mem[16'h1F59] = 8'hB5;
mem[16'h1F5A] = 8'hAC;
mem[16'h1F5B] = 8'hD4;
mem[16'h1F5C] = 8'hB5;
mem[16'h1F5D] = 8'h60;
mem[16'h1F5E] = 8'h08;
mem[16'h1F5F] = 8'h20;
mem[16'h1F60] = 8'h34;
mem[16'h1F61] = 8'hAF;
mem[16'h1F62] = 8'h20;
mem[16'h1F63] = 8'h4B;
mem[16'h1F64] = 8'hAF;
mem[16'h1F65] = 8'h20;
mem[16'h1F66] = 8'h0C;
mem[16'h1F67] = 8'hAF;
mem[16'h1F68] = 8'h28;
mem[16'h1F69] = 8'hB0;
mem[16'h1F6A] = 8'h09;
mem[16'h1F6B] = 8'hAE;
mem[16'h1F6C] = 8'hD1;
mem[16'h1F6D] = 8'hB5;
mem[16'h1F6E] = 8'hAC;
mem[16'h1F6F] = 8'hD2;
mem[16'h1F70] = 8'hB5;
mem[16'h1F71] = 8'h4C;
mem[16'h1F72] = 8'hB5;
mem[16'h1F73] = 8'hAF;
mem[16'h1F74] = 8'hA0;
mem[16'h1F75] = 8'h01;
mem[16'h1F76] = 8'hB1;
mem[16'h1F77] = 8'h42;
mem[16'h1F78] = 8'hF0;
mem[16'h1F79] = 8'h08;
mem[16'h1F7A] = 8'hAA;
mem[16'h1F7B] = 8'hC8;
mem[16'h1F7C] = 8'hB1;
mem[16'h1F7D] = 8'h42;
mem[16'h1F7E] = 8'hA8;
mem[16'h1F7F] = 8'h4C;
mem[16'h1F80] = 8'hB5;
mem[16'h1F81] = 8'hAF;
mem[16'h1F82] = 8'hAD;
mem[16'h1F83] = 8'hBB;
mem[16'h1F84] = 8'hB5;
mem[16'h1F85] = 8'hC9;
mem[16'h1F86] = 8'h04;
mem[16'h1F87] = 8'hF0;
mem[16'h1F88] = 8'h02;
mem[16'h1F89] = 8'h38;
mem[16'h1F8A] = 8'h60;
mem[16'h1F8B] = 8'h20;
mem[16'h1F8C] = 8'h44;
mem[16'h1F8D] = 8'hB2;
mem[16'h1F8E] = 8'hA0;
mem[16'h1F8F] = 8'h02;
mem[16'h1F90] = 8'h91;
mem[16'h1F91] = 8'h42;
mem[16'h1F92] = 8'h48;
mem[16'h1F93] = 8'h88;
mem[16'h1F94] = 8'hAD;
mem[16'h1F95] = 8'hF1;
mem[16'h1F96] = 8'hB5;
mem[16'h1F97] = 8'h91;
mem[16'h1F98] = 8'h42;
mem[16'h1F99] = 8'h48;
mem[16'h1F9A] = 8'h20;
mem[16'h1F9B] = 8'h3A;
mem[16'h1F9C] = 8'hAF;
mem[16'h1F9D] = 8'h20;
mem[16'h1F9E] = 8'hD6;
mem[16'h1F9F] = 8'hB7;
mem[16'h1FA0] = 8'hA0;
mem[16'h1FA1] = 8'h05;
mem[16'h1FA2] = 8'hAD;
mem[16'h1FA3] = 8'hDE;
mem[16'h1FA4] = 8'hB5;
mem[16'h1FA5] = 8'h91;
mem[16'h1FA6] = 8'h42;
mem[16'h1FA7] = 8'hC8;
mem[16'h1FA8] = 8'hAD;
mem[16'h1FA9] = 8'hDF;
mem[16'h1FAA] = 8'hB5;
mem[16'h1FAB] = 8'h91;
mem[16'h1FAC] = 8'h42;
mem[16'h1FAD] = 8'h68;
mem[16'h1FAE] = 8'hAA;
mem[16'h1FAF] = 8'h68;
mem[16'h1FB0] = 8'hA8;
mem[16'h1FB1] = 8'hA9;
mem[16'h1FB2] = 8'h02;
mem[16'h1FB3] = 8'hD0;
mem[16'h1FB4] = 8'h02;
mem[16'h1FB5] = 8'hA9;
mem[16'h1FB6] = 8'h01;
mem[16'h1FB7] = 8'h8E;
mem[16'h1FB8] = 8'hD3;
mem[16'h1FB9] = 8'hB5;
mem[16'h1FBA] = 8'h8C;
mem[16'h1FBB] = 8'hD4;
mem[16'h1FBC] = 8'hB5;
mem[16'h1FBD] = 8'h20;
mem[16'h1FBE] = 8'h52;
mem[16'h1FBF] = 8'hB0;
mem[16'h1FC0] = 8'hA0;
mem[16'h1FC1] = 8'h05;
mem[16'h1FC2] = 8'hB1;
mem[16'h1FC3] = 8'h42;
mem[16'h1FC4] = 8'h8D;
mem[16'h1FC5] = 8'hDC;
mem[16'h1FC6] = 8'hB5;
mem[16'h1FC7] = 8'h18;
mem[16'h1FC8] = 8'h6D;
mem[16'h1FC9] = 8'hDA;
mem[16'h1FCA] = 8'hB5;
mem[16'h1FCB] = 8'h8D;
mem[16'h1FCC] = 8'hDE;
mem[16'h1FCD] = 8'hB5;
mem[16'h1FCE] = 8'hC8;
mem[16'h1FCF] = 8'hB1;
mem[16'h1FD0] = 8'h42;
mem[16'h1FD1] = 8'h8D;
mem[16'h1FD2] = 8'hDD;
mem[16'h1FD3] = 8'hB5;
mem[16'h1FD4] = 8'h6D;
mem[16'h1FD5] = 8'hDB;
mem[16'h1FD6] = 8'hB5;
mem[16'h1FD7] = 8'h8D;
mem[16'h1FD8] = 8'hDF;
mem[16'h1FD9] = 8'hB5;
mem[16'h1FDA] = 8'h18;
mem[16'h1FDB] = 8'h60;
mem[16'h1FDC] = 8'h20;
mem[16'h1FDD] = 8'hE4;
mem[16'h1FDE] = 8'hAF;
mem[16'h1FDF] = 8'hA9;
mem[16'h1FE0] = 8'h01;
mem[16'h1FE1] = 8'h4C;
mem[16'h1FE2] = 8'h52;
mem[16'h1FE3] = 8'hB0;
mem[16'h1FE4] = 8'hAC;
mem[16'h1FE5] = 8'hCB;
mem[16'h1FE6] = 8'hB5;
mem[16'h1FE7] = 8'hAD;
mem[16'h1FE8] = 8'hCC;
mem[16'h1FE9] = 8'hB5;
mem[16'h1FEA] = 8'h8C;
mem[16'h1FEB] = 8'hF0;
mem[16'h1FEC] = 8'hB7;
mem[16'h1FED] = 8'h8D;
mem[16'h1FEE] = 8'hF1;
mem[16'h1FEF] = 8'hB7;
mem[16'h1FF0] = 8'hAE;
mem[16'h1FF1] = 8'hD6;
mem[16'h1FF2] = 8'hB5;
mem[16'h1FF3] = 8'hAC;
mem[16'h1FF4] = 8'hD7;
mem[16'h1FF5] = 8'hB5;
mem[16'h1FF6] = 8'h60;
mem[16'h1FF7] = 8'hA9;
mem[16'h1FF8] = 8'h01;
mem[16'h1FF9] = 8'hD0;
mem[16'h1FFA] = 8'h02;
mem[16'h1FFB] = 8'hA9;
mem[16'h1FFC] = 8'h02;
mem[16'h1FFD] = 8'hAC;
mem[16'h1FFE] = 8'hC3;
mem[16'h1FFF] = 8'hAA;
mem[16'h2000] = 8'h00;
mem[16'h2001] = 8'h42;
mem[16'h2002] = 8'h10;
mem[16'h2003] = 8'h00;
mem[16'h2004] = 8'h3C;
mem[16'h2005] = 8'h00;
mem[16'h2006] = 8'h00;
mem[16'h2007] = 8'h00;
mem[16'h2008] = 8'h00;
mem[16'h2009] = 8'h00;
mem[16'h200A] = 8'h3C;
mem[16'h200B] = 8'h3C;
mem[16'h200C] = 8'h3C;
mem[16'h200D] = 8'h3C;
mem[16'h200E] = 8'h3C;
mem[16'h200F] = 8'h3C;
mem[16'h2010] = 8'h00;
mem[16'h2011] = 8'h00;
mem[16'h2012] = 8'h00;
mem[16'h2013] = 8'h00;
mem[16'h2014] = 8'h44;
mem[16'h2015] = 8'h00;
mem[16'h2016] = 8'h00;
mem[16'h2017] = 8'h00;
mem[16'h2018] = 8'h00;
mem[16'h2019] = 8'h3C;
mem[16'h201A] = 8'h00;
mem[16'h201B] = 8'h00;
mem[16'h201C] = 8'h00;
mem[16'h201D] = 8'h00;
mem[16'h201E] = 8'h00;
mem[16'h201F] = 8'h3C;
mem[16'h2020] = 8'h3C;
mem[16'h2021] = 8'h3C;
mem[16'h2022] = 8'h3C;
mem[16'h2023] = 8'h3C;
mem[16'h2024] = 8'h3C;
mem[16'h2025] = 8'h00;
mem[16'h2026] = 8'h00;
mem[16'h2027] = 8'h00;
mem[16'h2028] = 8'hD5;
mem[16'h2029] = 8'hAA;
mem[16'h202A] = 8'hD5;
mem[16'h202B] = 8'hAA;
mem[16'h202C] = 8'hD5;
mem[16'h202D] = 8'hAA;
mem[16'h202E] = 8'hD5;
mem[16'h202F] = 8'hAA;
mem[16'h2030] = 8'hD5;
mem[16'h2031] = 8'hAA;
mem[16'h2032] = 8'hD5;
mem[16'h2033] = 8'hAA;
mem[16'h2034] = 8'hD5;
mem[16'h2035] = 8'hAA;
mem[16'h2036] = 8'hD5;
mem[16'h2037] = 8'hAA;
mem[16'h2038] = 8'hD5;
mem[16'h2039] = 8'hAA;
mem[16'h203A] = 8'hD5;
mem[16'h203B] = 8'hAA;
mem[16'h203C] = 8'hD5;
mem[16'h203D] = 8'hAA;
mem[16'h203E] = 8'hD5;
mem[16'h203F] = 8'hAA;
mem[16'h2040] = 8'hD5;
mem[16'h2041] = 8'hAA;
mem[16'h2042] = 8'hD5;
mem[16'h2043] = 8'hAA;
mem[16'h2044] = 8'hD5;
mem[16'h2045] = 8'hAA;
mem[16'h2046] = 8'hD5;
mem[16'h2047] = 8'hAA;
mem[16'h2048] = 8'hD5;
mem[16'h2049] = 8'hAA;
mem[16'h204A] = 8'hD5;
mem[16'h204B] = 8'hAA;
mem[16'h204C] = 8'h85;
mem[16'h204D] = 8'h00;
mem[16'h204E] = 8'h00;
mem[16'h204F] = 8'h00;
mem[16'h2050] = 8'h00;
mem[16'h2051] = 8'hF0;
mem[16'h2052] = 8'hC0;
mem[16'h2053] = 8'h83;
mem[16'h2054] = 8'h00;
mem[16'h2055] = 8'h00;
mem[16'h2056] = 8'h00;
mem[16'h2057] = 8'h00;
mem[16'h2058] = 8'h00;
mem[16'h2059] = 8'h00;
mem[16'h205A] = 8'h00;
mem[16'h205B] = 8'h00;
mem[16'h205C] = 8'h00;
mem[16'h205D] = 8'h00;
mem[16'h205E] = 8'h00;
mem[16'h205F] = 8'h00;
mem[16'h2060] = 8'h00;
mem[16'h2061] = 8'h00;
mem[16'h2062] = 8'h00;
mem[16'h2063] = 8'h00;
mem[16'h2064] = 8'h00;
mem[16'h2065] = 8'h00;
mem[16'h2066] = 8'h00;
mem[16'h2067] = 8'h00;
mem[16'h2068] = 8'h00;
mem[16'h2069] = 8'h00;
mem[16'h206A] = 8'h00;
mem[16'h206B] = 8'h00;
mem[16'h206C] = 8'h00;
mem[16'h206D] = 8'h00;
mem[16'h206E] = 8'h00;
mem[16'h206F] = 8'h00;
mem[16'h2070] = 8'h00;
mem[16'h2071] = 8'h00;
mem[16'h2072] = 8'h00;
mem[16'h2073] = 8'h00;
mem[16'h2074] = 8'h00;
mem[16'h2075] = 8'h00;
mem[16'h2076] = 8'h00;
mem[16'h2077] = 8'h2A;
mem[16'h2078] = 8'h00;
mem[16'h2079] = 8'h00;
mem[16'h207A] = 8'h00;
mem[16'h207B] = 8'h00;
mem[16'h207C] = 8'h00;
mem[16'h207D] = 8'h00;
mem[16'h207E] = 8'h00;
mem[16'h207F] = 8'h00;
mem[16'h2080] = 8'h02;
mem[16'h2081] = 8'h55;
mem[16'h2082] = 8'h28;
mem[16'h2083] = 8'h15;
mem[16'h2084] = 8'h2A;
mem[16'h2085] = 8'h11;
mem[16'h2086] = 8'h2A;
mem[16'h2087] = 8'h05;
mem[16'h2088] = 8'h02;
mem[16'h2089] = 8'h55;
mem[16'h208A] = 8'h28;
mem[16'h208B] = 8'h15;
mem[16'h208C] = 8'h2A;
mem[16'h208D] = 8'h11;
mem[16'h208E] = 8'h2A;
mem[16'h208F] = 8'h05;
mem[16'h2090] = 8'h02;
mem[16'h2091] = 8'h55;
mem[16'h2092] = 8'h28;
mem[16'h2093] = 8'h15;
mem[16'h2094] = 8'h2A;
mem[16'h2095] = 8'h11;
mem[16'h2096] = 8'h2A;
mem[16'h2097] = 8'h05;
mem[16'h2098] = 8'h02;
mem[16'h2099] = 8'h55;
mem[16'h209A] = 8'h28;
mem[16'h209B] = 8'h15;
mem[16'h209C] = 8'h2A;
mem[16'h209D] = 8'h11;
mem[16'h209E] = 8'h2A;
mem[16'h209F] = 8'h05;
mem[16'h20A0] = 8'h02;
mem[16'h20A1] = 8'h55;
mem[16'h20A2] = 8'h28;
mem[16'h20A3] = 8'h15;
mem[16'h20A4] = 8'h0A;
mem[16'h20A5] = 8'h00;
mem[16'h20A6] = 8'h70;
mem[16'h20A7] = 8'h07;
mem[16'h20A8] = 8'hD5;
mem[16'h20A9] = 8'hAA;
mem[16'h20AA] = 8'hD5;
mem[16'h20AB] = 8'hAA;
mem[16'h20AC] = 8'hD5;
mem[16'h20AD] = 8'hD5;
mem[16'h20AE] = 8'hAA;
mem[16'h20AF] = 8'hD5;
mem[16'h20B0] = 8'hAA;
mem[16'h20B1] = 8'hD5;
mem[16'h20B2] = 8'hAA;
mem[16'h20B3] = 8'hD5;
mem[16'h20B4] = 8'hD5;
mem[16'h20B5] = 8'hAA;
mem[16'h20B6] = 8'hD5;
mem[16'h20B7] = 8'hAA;
mem[16'h20B8] = 8'hD5;
mem[16'h20B9] = 8'hD6;
mem[16'h20BA] = 8'hAA;
mem[16'h20BB] = 8'hD5;
mem[16'h20BC] = 8'hAA;
mem[16'h20BD] = 8'hD5;
mem[16'h20BE] = 8'hAA;
mem[16'h20BF] = 8'hD5;
mem[16'h20C0] = 8'hD6;
mem[16'h20C1] = 8'hAA;
mem[16'h20C2] = 8'hD5;
mem[16'h20C3] = 8'hAA;
mem[16'h20C4] = 8'hAD;
mem[16'h20C5] = 8'hD5;
mem[16'h20C6] = 8'hAA;
mem[16'h20C7] = 8'hD5;
mem[16'h20C8] = 8'hAA;
mem[16'h20C9] = 8'hD5;
mem[16'h20CA] = 8'hAA;
mem[16'h20CB] = 8'hAD;
mem[16'h20CC] = 8'h85;
mem[16'h20CD] = 8'h00;
mem[16'h20CE] = 8'h00;
mem[16'h20CF] = 8'h2A;
mem[16'h20D0] = 8'h00;
mem[16'h20D1] = 8'h00;
mem[16'h20D2] = 8'h00;
mem[16'h20D3] = 8'h00;
mem[16'h20D4] = 8'h00;
mem[16'h20D5] = 8'h54;
mem[16'h20D6] = 8'h2A;
mem[16'h20D7] = 8'h03;
mem[16'h20D8] = 8'h00;
mem[16'h20D9] = 8'h00;
mem[16'h20DA] = 8'h00;
mem[16'h20DB] = 8'h00;
mem[16'h20DC] = 8'h00;
mem[16'h20DD] = 8'h00;
mem[16'h20DE] = 8'h00;
mem[16'h20DF] = 8'h00;
mem[16'h20E0] = 8'h00;
mem[16'h20E1] = 8'h54;
mem[16'h20E2] = 8'h2A;
mem[16'h20E3] = 8'h03;
mem[16'h20E4] = 8'h00;
mem[16'h20E5] = 8'h00;
mem[16'h20E6] = 8'h00;
mem[16'h20E7] = 8'h00;
mem[16'h20E8] = 8'h00;
mem[16'h20E9] = 8'h00;
mem[16'h20EA] = 8'h00;
mem[16'h20EB] = 8'h00;
mem[16'h20EC] = 8'h00;
mem[16'h20ED] = 8'h54;
mem[16'h20EE] = 8'h2A;
mem[16'h20EF] = 8'h03;
mem[16'h20F0] = 8'h00;
mem[16'h20F1] = 8'h00;
mem[16'h20F2] = 8'h00;
mem[16'h20F3] = 8'h00;
mem[16'h20F4] = 8'h00;
mem[16'h20F5] = 8'h00;
mem[16'h20F6] = 8'h00;
mem[16'h20F7] = 8'h2A;
mem[16'h20F8] = 8'h00;
mem[16'h20F9] = 8'h00;
mem[16'h20FA] = 8'h00;
mem[16'h20FB] = 8'h00;
mem[16'h20FC] = 8'h00;
mem[16'h20FD] = 8'h00;
mem[16'h20FE] = 8'h00;
mem[16'h20FF] = 8'h00;
mem[16'h2100] = 8'h2A;
mem[16'h2101] = 8'h45;
mem[16'h2102] = 8'h2A;
mem[16'h2103] = 8'hAA;
mem[16'h2104] = 8'hD5;
mem[16'h2105] = 8'h41;
mem[16'h2106] = 8'h20;
mem[16'h2107] = 8'h15;
mem[16'h2108] = 8'h2A;
mem[16'h2109] = 8'h45;
mem[16'h210A] = 8'hD5;
mem[16'h210B] = 8'hAA;
mem[16'h210C] = 8'h2A;
mem[16'h210D] = 8'h41;
mem[16'h210E] = 8'h20;
mem[16'h210F] = 8'h15;
mem[16'h2110] = 8'hD5;
mem[16'h2111] = 8'hAA;
mem[16'h2112] = 8'h2A;
mem[16'h2113] = 8'h44;
mem[16'h2114] = 8'h2A;
mem[16'h2115] = 8'h41;
mem[16'h2116] = 8'h20;
mem[16'h2117] = 8'hAA;
mem[16'h2118] = 8'hD5;
mem[16'h2119] = 8'h45;
mem[16'h211A] = 8'h2A;
mem[16'h211B] = 8'h44;
mem[16'h211C] = 8'h2A;
mem[16'h211D] = 8'hAA;
mem[16'h211E] = 8'hD5;
mem[16'h211F] = 8'h15;
mem[16'h2120] = 8'h2A;
mem[16'h2121] = 8'h45;
mem[16'h2122] = 8'h2A;
mem[16'h2123] = 8'h44;
mem[16'h2124] = 8'h0A;
mem[16'h2125] = 8'h00;
mem[16'h2126] = 8'h00;
mem[16'h2127] = 8'h00;
mem[16'h2128] = 8'hD5;
mem[16'h2129] = 8'hAA;
mem[16'h212A] = 8'hD5;
mem[16'h212B] = 8'hAA;
mem[16'h212C] = 8'hD5;
mem[16'h212D] = 8'hCF;
mem[16'h212E] = 8'hAA;
mem[16'h212F] = 8'hFA;
mem[16'h2130] = 8'hA9;
mem[16'h2131] = 8'hA5;
mem[16'h2132] = 8'h9F;
mem[16'h2133] = 8'hD5;
mem[16'h2134] = 8'hD4;
mem[16'h2135] = 8'hAA;
mem[16'h2136] = 8'hD5;
mem[16'h2137] = 8'hAA;
mem[16'h2138] = 8'hD5;
mem[16'h2139] = 8'hAA;
mem[16'h213A] = 8'hD5;
mem[16'h213B] = 8'hEA;
mem[16'h213C] = 8'hA7;
mem[16'h213D] = 8'h95;
mem[16'h213E] = 8'hFD;
mem[16'h213F] = 8'hD4;
mem[16'h2140] = 8'hD2;
mem[16'h2141] = 8'hCF;
mem[16'h2142] = 8'hAA;
mem[16'h2143] = 8'hAA;
mem[16'h2144] = 8'hD5;
mem[16'h2145] = 8'hAA;
mem[16'h2146] = 8'hD5;
mem[16'h2147] = 8'hAA;
mem[16'h2148] = 8'hD5;
mem[16'h2149] = 8'hAA;
mem[16'h214A] = 8'hD5;
mem[16'h214B] = 8'hAA;
mem[16'h214C] = 8'h85;
mem[16'h214D] = 8'h00;
mem[16'h214E] = 8'h00;
mem[16'h214F] = 8'h2A;
mem[16'h2150] = 8'h00;
mem[16'h2151] = 8'h00;
mem[16'h2152] = 8'h00;
mem[16'h2153] = 8'h00;
mem[16'h2154] = 8'h00;
mem[16'h2155] = 8'h00;
mem[16'h2156] = 8'h00;
mem[16'h2157] = 8'h00;
mem[16'h2158] = 8'h00;
mem[16'h2159] = 8'h00;
mem[16'h215A] = 8'h00;
mem[16'h215B] = 8'h00;
mem[16'h215C] = 8'h00;
mem[16'h215D] = 8'h00;
mem[16'h215E] = 8'h00;
mem[16'h215F] = 8'h00;
mem[16'h2160] = 8'h00;
mem[16'h2161] = 8'h00;
mem[16'h2162] = 8'h00;
mem[16'h2163] = 8'h00;
mem[16'h2164] = 8'h00;
mem[16'h2165] = 8'h00;
mem[16'h2166] = 8'h00;
mem[16'h2167] = 8'h00;
mem[16'h2168] = 8'h00;
mem[16'h2169] = 8'h00;
mem[16'h216A] = 8'h00;
mem[16'h216B] = 8'h00;
mem[16'h216C] = 8'h00;
mem[16'h216D] = 8'h00;
mem[16'h216E] = 8'h00;
mem[16'h216F] = 8'h00;
mem[16'h2170] = 8'h00;
mem[16'h2171] = 8'h00;
mem[16'h2172] = 8'h00;
mem[16'h2173] = 8'h00;
mem[16'h2174] = 8'h00;
mem[16'h2175] = 8'h00;
mem[16'h2176] = 8'h00;
mem[16'h2177] = 8'h2A;
mem[16'h2178] = 8'h00;
mem[16'h2179] = 8'h00;
mem[16'h217A] = 8'h00;
mem[16'h217B] = 8'h00;
mem[16'h217C] = 8'h00;
mem[16'h217D] = 8'h00;
mem[16'h217E] = 8'h00;
mem[16'h217F] = 8'h00;
mem[16'h2180] = 8'hD5;
mem[16'h2181] = 8'hAA;
mem[16'h2182] = 8'hD5;
mem[16'h2183] = 8'hAA;
mem[16'h2184] = 8'hD5;
mem[16'h2185] = 8'hAA;
mem[16'h2186] = 8'hAD;
mem[16'h2187] = 8'hD5;
mem[16'h2188] = 8'hAA;
mem[16'h2189] = 8'hD5;
mem[16'h218A] = 8'hAA;
mem[16'h218B] = 8'hD5;
mem[16'h218C] = 8'hAA;
mem[16'h218D] = 8'hD5;
mem[16'h218E] = 8'hAA;
mem[16'h218F] = 8'hB5;
mem[16'h2190] = 8'hD5;
mem[16'h2191] = 8'hAA;
mem[16'h2192] = 8'hB5;
mem[16'h2193] = 8'hD5;
mem[16'h2194] = 8'hAA;
mem[16'h2195] = 8'hD5;
mem[16'h2196] = 8'hAA;
mem[16'h2197] = 8'hD5;
mem[16'h2198] = 8'hAA;
mem[16'h2199] = 8'hD5;
mem[16'h219A] = 8'hAA;
mem[16'h219B] = 8'hD5;
mem[16'h219C] = 8'hD5;
mem[16'h219D] = 8'hAA;
mem[16'h219E] = 8'hD5;
mem[16'h219F] = 8'hAA;
mem[16'h21A0] = 8'hD5;
mem[16'h21A1] = 8'hAA;
mem[16'h21A2] = 8'hD5;
mem[16'h21A3] = 8'hAA;
mem[16'h21A4] = 8'h85;
mem[16'h21A5] = 8'h00;
mem[16'h21A6] = 8'h7C;
mem[16'h21A7] = 8'h1F;
mem[16'h21A8] = 8'hD5;
mem[16'h21A9] = 8'hAA;
mem[16'h21AA] = 8'hD5;
mem[16'h21AB] = 8'hAA;
mem[16'h21AC] = 8'hD5;
mem[16'h21AD] = 8'hAA;
mem[16'h21AE] = 8'hD5;
mem[16'h21AF] = 8'hAA;
mem[16'h21B0] = 8'hD5;
mem[16'h21B1] = 8'hAA;
mem[16'h21B2] = 8'hD5;
mem[16'h21B3] = 8'hAA;
mem[16'h21B4] = 8'hD5;
mem[16'h21B5] = 8'hAA;
mem[16'h21B6] = 8'hD5;
mem[16'h21B7] = 8'hAA;
mem[16'h21B8] = 8'hD5;
mem[16'h21B9] = 8'hAA;
mem[16'h21BA] = 8'hD5;
mem[16'h21BB] = 8'hAA;
mem[16'h21BC] = 8'hD5;
mem[16'h21BD] = 8'hAA;
mem[16'h21BE] = 8'hD5;
mem[16'h21BF] = 8'hAA;
mem[16'h21C0] = 8'hD5;
mem[16'h21C1] = 8'hAA;
mem[16'h21C2] = 8'hD5;
mem[16'h21C3] = 8'hAA;
mem[16'h21C4] = 8'hD5;
mem[16'h21C5] = 8'hAA;
mem[16'h21C6] = 8'hD5;
mem[16'h21C7] = 8'hAA;
mem[16'h21C8] = 8'hD5;
mem[16'h21C9] = 8'hAA;
mem[16'h21CA] = 8'hD5;
mem[16'h21CB] = 8'hAA;
mem[16'h21CC] = 8'h85;
mem[16'h21CD] = 8'h00;
mem[16'h21CE] = 8'h00;
mem[16'h21CF] = 8'h2A;
mem[16'h21D0] = 8'h00;
mem[16'h21D1] = 8'hA8;
mem[16'h21D2] = 8'hF5;
mem[16'h21D3] = 8'h81;
mem[16'h21D4] = 8'h00;
mem[16'h21D5] = 8'h00;
mem[16'h21D6] = 8'h00;
mem[16'h21D7] = 8'h00;
mem[16'h21D8] = 8'h00;
mem[16'h21D9] = 8'h00;
mem[16'h21DA] = 8'h00;
mem[16'h21DB] = 8'hC0;
mem[16'h21DC] = 8'hAA;
mem[16'h21DD] = 8'h8F;
mem[16'h21DE] = 8'h00;
mem[16'h21DF] = 8'h00;
mem[16'h21E0] = 8'h00;
mem[16'h21E1] = 8'h00;
mem[16'h21E2] = 8'h00;
mem[16'h21E3] = 8'h00;
mem[16'h21E4] = 8'h00;
mem[16'h21E5] = 8'h00;
mem[16'h21E6] = 8'hD4;
mem[16'h21E7] = 8'hFA;
mem[16'h21E8] = 8'h80;
mem[16'h21E9] = 8'h00;
mem[16'h21EA] = 8'h00;
mem[16'h21EB] = 8'h00;
mem[16'h21EC] = 8'h00;
mem[16'h21ED] = 8'h00;
mem[16'h21EE] = 8'h00;
mem[16'h21EF] = 8'h00;
mem[16'h21F0] = 8'h00;
mem[16'h21F1] = 8'h00;
mem[16'h21F2] = 8'h00;
mem[16'h21F3] = 8'h00;
mem[16'h21F4] = 8'h00;
mem[16'h21F5] = 8'h00;
mem[16'h21F6] = 8'h00;
mem[16'h21F7] = 8'h2A;
mem[16'h21F8] = 8'h00;
mem[16'h21F9] = 8'h00;
mem[16'h21FA] = 8'h00;
mem[16'h21FB] = 8'h00;
mem[16'h21FC] = 8'h00;
mem[16'h21FD] = 8'h00;
mem[16'h21FE] = 8'h00;
mem[16'h21FF] = 8'h00;
mem[16'h2200] = 8'hD5;
mem[16'h2201] = 8'hAA;
mem[16'h2202] = 8'hD5;
mem[16'h2203] = 8'hAA;
mem[16'h2204] = 8'hD5;
mem[16'h2205] = 8'hAA;
mem[16'h2206] = 8'hD5;
mem[16'h2207] = 8'hAA;
mem[16'h2208] = 8'hD5;
mem[16'h2209] = 8'hAA;
mem[16'h220A] = 8'hD5;
mem[16'h220B] = 8'hAA;
mem[16'h220C] = 8'hD5;
mem[16'h220D] = 8'hAA;
mem[16'h220E] = 8'hD5;
mem[16'h220F] = 8'hAA;
mem[16'h2210] = 8'hD5;
mem[16'h2211] = 8'hAA;
mem[16'h2212] = 8'hD5;
mem[16'h2213] = 8'hAA;
mem[16'h2214] = 8'hD5;
mem[16'h2215] = 8'hAA;
mem[16'h2216] = 8'hD5;
mem[16'h2217] = 8'hAA;
mem[16'h2218] = 8'hD5;
mem[16'h2219] = 8'hAA;
mem[16'h221A] = 8'hD5;
mem[16'h221B] = 8'hAA;
mem[16'h221C] = 8'hD5;
mem[16'h221D] = 8'hAA;
mem[16'h221E] = 8'hD5;
mem[16'h221F] = 8'hAA;
mem[16'h2220] = 8'hD5;
mem[16'h2221] = 8'hAA;
mem[16'h2222] = 8'hD5;
mem[16'h2223] = 8'hAA;
mem[16'h2224] = 8'h85;
mem[16'h2225] = 8'h00;
mem[16'h2226] = 8'h60;
mem[16'h2227] = 8'h03;
mem[16'h2228] = 8'h22;
mem[16'h2229] = 8'h15;
mem[16'h222A] = 8'h22;
mem[16'h222B] = 8'h55;
mem[16'h222C] = 8'h20;
mem[16'h222D] = 8'h50;
mem[16'h222E] = 8'h0A;
mem[16'h222F] = 8'h55;
mem[16'h2230] = 8'h22;
mem[16'h2231] = 8'h15;
mem[16'h2232] = 8'h22;
mem[16'h2233] = 8'h55;
mem[16'h2234] = 8'h20;
mem[16'h2235] = 8'h50;
mem[16'h2236] = 8'h0A;
mem[16'h2237] = 8'h55;
mem[16'h2238] = 8'h22;
mem[16'h2239] = 8'h15;
mem[16'h223A] = 8'h22;
mem[16'h223B] = 8'h55;
mem[16'h223C] = 8'h20;
mem[16'h223D] = 8'h50;
mem[16'h223E] = 8'h0A;
mem[16'h223F] = 8'h55;
mem[16'h2240] = 8'h22;
mem[16'h2241] = 8'h15;
mem[16'h2242] = 8'h22;
mem[16'h2243] = 8'h55;
mem[16'h2244] = 8'h20;
mem[16'h2245] = 8'h50;
mem[16'h2246] = 8'h0A;
mem[16'h2247] = 8'h55;
mem[16'h2248] = 8'h22;
mem[16'h2249] = 8'h15;
mem[16'h224A] = 8'h22;
mem[16'h224B] = 8'h55;
mem[16'h224C] = 8'h00;
mem[16'h224D] = 8'h00;
mem[16'h224E] = 8'h00;
mem[16'h224F] = 8'h2A;
mem[16'h2250] = 8'h00;
mem[16'h2251] = 8'h00;
mem[16'h2252] = 8'h00;
mem[16'h2253] = 8'h00;
mem[16'h2254] = 8'h00;
mem[16'h2255] = 8'h00;
mem[16'h2256] = 8'h00;
mem[16'h2257] = 8'h00;
mem[16'h2258] = 8'h00;
mem[16'h2259] = 8'h00;
mem[16'h225A] = 8'h00;
mem[16'h225B] = 8'h00;
mem[16'h225C] = 8'h00;
mem[16'h225D] = 8'h00;
mem[16'h225E] = 8'h00;
mem[16'h225F] = 8'h00;
mem[16'h2260] = 8'h00;
mem[16'h2261] = 8'h00;
mem[16'h2262] = 8'h00;
mem[16'h2263] = 8'h00;
mem[16'h2264] = 8'h00;
mem[16'h2265] = 8'h00;
mem[16'h2266] = 8'h00;
mem[16'h2267] = 8'h00;
mem[16'h2268] = 8'h00;
mem[16'h2269] = 8'h00;
mem[16'h226A] = 8'h00;
mem[16'h226B] = 8'h00;
mem[16'h226C] = 8'h00;
mem[16'h226D] = 8'h00;
mem[16'h226E] = 8'h00;
mem[16'h226F] = 8'h00;
mem[16'h2270] = 8'h00;
mem[16'h2271] = 8'h00;
mem[16'h2272] = 8'h00;
mem[16'h2273] = 8'h00;
mem[16'h2274] = 8'h00;
mem[16'h2275] = 8'h00;
mem[16'h2276] = 8'h00;
mem[16'h2277] = 8'h2A;
mem[16'h2278] = 8'h00;
mem[16'h2279] = 8'h00;
mem[16'h227A] = 8'h00;
mem[16'h227B] = 8'h00;
mem[16'h227C] = 8'h00;
mem[16'h227D] = 8'h00;
mem[16'h227E] = 8'h00;
mem[16'h227F] = 8'h00;
mem[16'h2280] = 8'hB5;
mem[16'h2281] = 8'hD5;
mem[16'h2282] = 8'hD4;
mem[16'h2283] = 8'hD6;
mem[16'h2284] = 8'hCA;
mem[16'h2285] = 8'hAA;
mem[16'h2286] = 8'hD5;
mem[16'h2287] = 8'hAA;
mem[16'h2288] = 8'hD5;
mem[16'h2289] = 8'hD5;
mem[16'h228A] = 8'hD2;
mem[16'h228B] = 8'hDA;
mem[16'h228C] = 8'hAA;
mem[16'h228D] = 8'hAA;
mem[16'h228E] = 8'hD5;
mem[16'h228F] = 8'hAA;
mem[16'h2290] = 8'hD5;
mem[16'h2291] = 8'hD6;
mem[16'h2292] = 8'hCA;
mem[16'h2293] = 8'hEA;
mem[16'h2294] = 8'hAA;
mem[16'h2295] = 8'hA9;
mem[16'h2296] = 8'hD5;
mem[16'h2297] = 8'hAA;
mem[16'h2298] = 8'hD5;
mem[16'h2299] = 8'hDA;
mem[16'h229A] = 8'hAA;
mem[16'h229B] = 8'hAA;
mem[16'h229C] = 8'hAB;
mem[16'h229D] = 8'hA5;
mem[16'h229E] = 8'hD5;
mem[16'h229F] = 8'hAA;
mem[16'h22A0] = 8'hD5;
mem[16'h22A1] = 8'hAA;
mem[16'h22A2] = 8'hD5;
mem[16'h22A3] = 8'hAA;
mem[16'h22A4] = 8'h85;
mem[16'h22A5] = 8'h00;
mem[16'h22A6] = 8'h44;
mem[16'h22A7] = 8'h12;
mem[16'h22A8] = 8'h28;
mem[16'h22A9] = 8'h15;
mem[16'h22AA] = 8'h08;
mem[16'h22AB] = 8'h54;
mem[16'h22AC] = 8'h22;
mem[16'h22AD] = 8'h55;
mem[16'h22AE] = 8'h28;
mem[16'h22AF] = 8'h45;
mem[16'h22B0] = 8'h28;
mem[16'h22B1] = 8'h15;
mem[16'h22B2] = 8'h08;
mem[16'h22B3] = 8'h54;
mem[16'h22B4] = 8'h22;
mem[16'h22B5] = 8'h55;
mem[16'h22B6] = 8'h28;
mem[16'h22B7] = 8'h45;
mem[16'h22B8] = 8'h28;
mem[16'h22B9] = 8'h15;
mem[16'h22BA] = 8'h08;
mem[16'h22BB] = 8'h54;
mem[16'h22BC] = 8'h22;
mem[16'h22BD] = 8'h55;
mem[16'h22BE] = 8'h28;
mem[16'h22BF] = 8'h45;
mem[16'h22C0] = 8'h28;
mem[16'h22C1] = 8'h15;
mem[16'h22C2] = 8'h08;
mem[16'h22C3] = 8'h54;
mem[16'h22C4] = 8'h22;
mem[16'h22C5] = 8'h55;
mem[16'h22C6] = 8'h28;
mem[16'h22C7] = 8'h45;
mem[16'h22C8] = 8'h28;
mem[16'h22C9] = 8'h15;
mem[16'h22CA] = 8'h08;
mem[16'h22CB] = 8'h54;
mem[16'h22CC] = 8'h02;
mem[16'h22CD] = 8'h00;
mem[16'h22CE] = 8'h00;
mem[16'h22CF] = 8'h2A;
mem[16'h22D0] = 8'h00;
mem[16'h22D1] = 8'h00;
mem[16'h22D2] = 8'h00;
mem[16'h22D3] = 8'h00;
mem[16'h22D4] = 8'h15;
mem[16'h22D5] = 8'h28;
mem[16'h22D6] = 8'h1D;
mem[16'h22D7] = 8'h00;
mem[16'h22D8] = 8'h00;
mem[16'h22D9] = 8'h00;
mem[16'h22DA] = 8'h00;
mem[16'h22DB] = 8'h00;
mem[16'h22DC] = 8'h00;
mem[16'h22DD] = 8'h00;
mem[16'h22DE] = 8'h00;
mem[16'h22DF] = 8'h00;
mem[16'h22E0] = 8'h00;
mem[16'h22E1] = 8'h00;
mem[16'h22E2] = 8'h15;
mem[16'h22E3] = 8'h28;
mem[16'h22E4] = 8'h1D;
mem[16'h22E5] = 8'h00;
mem[16'h22E6] = 8'h00;
mem[16'h22E7] = 8'h00;
mem[16'h22E8] = 8'h00;
mem[16'h22E9] = 8'h00;
mem[16'h22EA] = 8'h00;
mem[16'h22EB] = 8'h00;
mem[16'h22EC] = 8'h00;
mem[16'h22ED] = 8'h00;
mem[16'h22EE] = 8'h00;
mem[16'h22EF] = 8'h00;
mem[16'h22F0] = 8'h15;
mem[16'h22F1] = 8'h28;
mem[16'h22F2] = 8'h1D;
mem[16'h22F3] = 8'h00;
mem[16'h22F4] = 8'h00;
mem[16'h22F5] = 8'h00;
mem[16'h22F6] = 8'h00;
mem[16'h22F7] = 8'h2A;
mem[16'h22F8] = 8'h00;
mem[16'h22F9] = 8'h00;
mem[16'h22FA] = 8'h00;
mem[16'h22FB] = 8'h00;
mem[16'h22FC] = 8'h00;
mem[16'h22FD] = 8'h00;
mem[16'h22FE] = 8'h00;
mem[16'h22FF] = 8'h00;
mem[16'h2300] = 8'hD5;
mem[16'h2301] = 8'hAA;
mem[16'h2302] = 8'hD5;
mem[16'h2303] = 8'hAA;
mem[16'h2304] = 8'hD5;
mem[16'h2305] = 8'hAA;
mem[16'h2306] = 8'hD5;
mem[16'h2307] = 8'hAA;
mem[16'h2308] = 8'hD5;
mem[16'h2309] = 8'hAA;
mem[16'h230A] = 8'hD5;
mem[16'h230B] = 8'hAA;
mem[16'h230C] = 8'hD5;
mem[16'h230D] = 8'hAA;
mem[16'h230E] = 8'hD5;
mem[16'h230F] = 8'hAA;
mem[16'h2310] = 8'hD5;
mem[16'h2311] = 8'hAA;
mem[16'h2312] = 8'hD5;
mem[16'h2313] = 8'hAA;
mem[16'h2314] = 8'hD5;
mem[16'h2315] = 8'hAA;
mem[16'h2316] = 8'hD5;
mem[16'h2317] = 8'hAA;
mem[16'h2318] = 8'hD5;
mem[16'h2319] = 8'hAA;
mem[16'h231A] = 8'hD5;
mem[16'h231B] = 8'hAA;
mem[16'h231C] = 8'hD5;
mem[16'h231D] = 8'hAA;
mem[16'h231E] = 8'hD5;
mem[16'h231F] = 8'hAA;
mem[16'h2320] = 8'hD5;
mem[16'h2321] = 8'hAA;
mem[16'h2322] = 8'hD5;
mem[16'h2323] = 8'hAA;
mem[16'h2324] = 8'h85;
mem[16'h2325] = 8'h00;
mem[16'h2326] = 8'h40;
mem[16'h2327] = 8'h01;
mem[16'h2328] = 8'h00;
mem[16'h2329] = 8'h00;
mem[16'h232A] = 8'h7D;
mem[16'h232B] = 8'h55;
mem[16'h232C] = 8'h0A;
mem[16'h232D] = 8'h00;
mem[16'h232E] = 8'h00;
mem[16'h232F] = 8'h00;
mem[16'h2330] = 8'h00;
mem[16'h2331] = 8'h00;
mem[16'h2332] = 8'h00;
mem[16'h2333] = 8'h00;
mem[16'h2334] = 8'h00;
mem[16'h2335] = 8'h00;
mem[16'h2336] = 8'h00;
mem[16'h2337] = 8'h00;
mem[16'h2338] = 8'h7D;
mem[16'h2339] = 8'h55;
mem[16'h233A] = 8'h0A;
mem[16'h233B] = 8'h00;
mem[16'h233C] = 8'h00;
mem[16'h233D] = 8'h00;
mem[16'h233E] = 8'h00;
mem[16'h233F] = 8'h00;
mem[16'h2340] = 8'h00;
mem[16'h2341] = 8'h00;
mem[16'h2342] = 8'h00;
mem[16'h2343] = 8'h00;
mem[16'h2344] = 8'h00;
mem[16'h2345] = 8'h00;
mem[16'h2346] = 8'h00;
mem[16'h2347] = 8'h00;
mem[16'h2348] = 8'h00;
mem[16'h2349] = 8'h00;
mem[16'h234A] = 8'h00;
mem[16'h234B] = 8'h00;
mem[16'h234C] = 8'h00;
mem[16'h234D] = 8'h00;
mem[16'h234E] = 8'h00;
mem[16'h234F] = 8'h2A;
mem[16'h2350] = 8'h2A;
mem[16'h2351] = 8'h54;
mem[16'h2352] = 8'h0A;
mem[16'h2353] = 8'h55;
mem[16'h2354] = 8'h08;
mem[16'h2355] = 8'h55;
mem[16'h2356] = 8'h02;
mem[16'h2357] = 8'h41;
mem[16'h2358] = 8'h2A;
mem[16'h2359] = 8'h54;
mem[16'h235A] = 8'h0A;
mem[16'h235B] = 8'h55;
mem[16'h235C] = 8'h08;
mem[16'h235D] = 8'h55;
mem[16'h235E] = 8'h02;
mem[16'h235F] = 8'h41;
mem[16'h2360] = 8'h2A;
mem[16'h2361] = 8'h54;
mem[16'h2362] = 8'h40;
mem[16'h2363] = 8'h01;
mem[16'h2364] = 8'h08;
mem[16'h2365] = 8'h55;
mem[16'h2366] = 8'h02;
mem[16'h2367] = 8'h41;
mem[16'h2368] = 8'h2A;
mem[16'h2369] = 8'h54;
mem[16'h236A] = 8'h0A;
mem[16'h236B] = 8'h55;
mem[16'h236C] = 8'h08;
mem[16'h236D] = 8'h55;
mem[16'h236E] = 8'h02;
mem[16'h236F] = 8'h41;
mem[16'h2370] = 8'h2A;
mem[16'h2371] = 8'h54;
mem[16'h2372] = 8'h0A;
mem[16'h2373] = 8'h55;
mem[16'h2374] = 8'h08;
mem[16'h2375] = 8'h00;
mem[16'h2376] = 8'h00;
mem[16'h2377] = 8'h2A;
mem[16'h2378] = 8'h00;
mem[16'h2379] = 8'h00;
mem[16'h237A] = 8'h00;
mem[16'h237B] = 8'h00;
mem[16'h237C] = 8'h00;
mem[16'h237D] = 8'h00;
mem[16'h237E] = 8'h00;
mem[16'h237F] = 8'h00;
mem[16'h2380] = 8'hAB;
mem[16'h2381] = 8'hAD;
mem[16'h2382] = 8'hD5;
mem[16'h2383] = 8'hAA;
mem[16'h2384] = 8'hD5;
mem[16'h2385] = 8'hAA;
mem[16'h2386] = 8'hD5;
mem[16'h2387] = 8'hAA;
mem[16'h2388] = 8'hD5;
mem[16'h2389] = 8'hAA;
mem[16'h238A] = 8'hD5;
mem[16'h238B] = 8'hD5;
mem[16'h238C] = 8'hAA;
mem[16'h238D] = 8'hD5;
mem[16'h238E] = 8'hAA;
mem[16'h238F] = 8'hD5;
mem[16'h2390] = 8'hAA;
mem[16'h2391] = 8'hD5;
mem[16'h2392] = 8'hAA;
mem[16'h2393] = 8'hD5;
mem[16'h2394] = 8'hAA;
mem[16'h2395] = 8'hD5;
mem[16'h2396] = 8'hAA;
mem[16'h2397] = 8'hD5;
mem[16'h2398] = 8'hAA;
mem[16'h2399] = 8'hD5;
mem[16'h239A] = 8'hD5;
mem[16'h239B] = 8'hAA;
mem[16'h239C] = 8'hD5;
mem[16'h239D] = 8'hAA;
mem[16'h239E] = 8'hD5;
mem[16'h239F] = 8'hAA;
mem[16'h23A0] = 8'hD5;
mem[16'h23A1] = 8'hAA;
mem[16'h23A2] = 8'hD5;
mem[16'h23A3] = 8'hAA;
mem[16'h23A4] = 8'h85;
mem[16'h23A5] = 8'h00;
mem[16'h23A6] = 8'h0E;
mem[16'h23A7] = 8'h38;
mem[16'h23A8] = 8'h00;
mem[16'h23A9] = 8'h00;
mem[16'h23AA] = 8'h00;
mem[16'h23AB] = 8'h00;
mem[16'h23AC] = 8'h00;
mem[16'h23AD] = 8'h00;
mem[16'h23AE] = 8'h00;
mem[16'h23AF] = 8'h00;
mem[16'h23B0] = 8'h00;
mem[16'h23B1] = 8'h00;
mem[16'h23B2] = 8'h00;
mem[16'h23B3] = 8'h00;
mem[16'h23B4] = 8'h00;
mem[16'h23B5] = 8'h00;
mem[16'h23B6] = 8'h00;
mem[16'h23B7] = 8'h00;
mem[16'h23B8] = 8'h00;
mem[16'h23B9] = 8'h00;
mem[16'h23BA] = 8'h00;
mem[16'h23BB] = 8'h00;
mem[16'h23BC] = 8'h00;
mem[16'h23BD] = 8'h00;
mem[16'h23BE] = 8'h00;
mem[16'h23BF] = 8'h00;
mem[16'h23C0] = 8'h00;
mem[16'h23C1] = 8'h00;
mem[16'h23C2] = 8'h00;
mem[16'h23C3] = 8'h00;
mem[16'h23C4] = 8'h00;
mem[16'h23C5] = 8'h00;
mem[16'h23C6] = 8'h00;
mem[16'h23C7] = 8'h00;
mem[16'h23C8] = 8'h00;
mem[16'h23C9] = 8'h00;
mem[16'h23CA] = 8'h00;
mem[16'h23CB] = 8'h00;
mem[16'h23CC] = 8'h00;
mem[16'h23CD] = 8'h00;
mem[16'h23CE] = 8'h00;
mem[16'h23CF] = 8'h2A;
mem[16'h23D0] = 8'h22;
mem[16'h23D1] = 8'h15;
mem[16'h23D2] = 8'h22;
mem[16'h23D3] = 8'h55;
mem[16'h23D4] = 8'h20;
mem[16'h23D5] = 8'h50;
mem[16'h23D6] = 8'h0A;
mem[16'h23D7] = 8'h55;
mem[16'h23D8] = 8'h22;
mem[16'h23D9] = 8'h15;
mem[16'h23DA] = 8'h22;
mem[16'h23DB] = 8'h55;
mem[16'h23DC] = 8'h20;
mem[16'h23DD] = 8'h50;
mem[16'h23DE] = 8'h0A;
mem[16'h23DF] = 8'h55;
mem[16'h23E0] = 8'h22;
mem[16'h23E1] = 8'h15;
mem[16'h23E2] = 8'h7C;
mem[16'h23E3] = 8'h1F;
mem[16'h23E4] = 8'h20;
mem[16'h23E5] = 8'h50;
mem[16'h23E6] = 8'h0A;
mem[16'h23E7] = 8'h55;
mem[16'h23E8] = 8'h22;
mem[16'h23E9] = 8'h15;
mem[16'h23EA] = 8'h22;
mem[16'h23EB] = 8'h55;
mem[16'h23EC] = 8'h20;
mem[16'h23ED] = 8'h50;
mem[16'h23EE] = 8'h0A;
mem[16'h23EF] = 8'h55;
mem[16'h23F0] = 8'h22;
mem[16'h23F1] = 8'h15;
mem[16'h23F2] = 8'h22;
mem[16'h23F3] = 8'h55;
mem[16'h23F4] = 8'h00;
mem[16'h23F5] = 8'h42;
mem[16'h23F6] = 8'h00;
mem[16'h23F7] = 8'h2A;
mem[16'h23F8] = 8'h00;
mem[16'h23F9] = 8'h00;
mem[16'h23FA] = 8'h00;
mem[16'h23FB] = 8'h00;
mem[16'h23FC] = 8'h00;
mem[16'h23FD] = 8'h00;
mem[16'h23FE] = 8'h00;
mem[16'h23FF] = 8'h00;
mem[16'h2400] = 8'h00;
mem[16'h2401] = 8'h42;
mem[16'h2402] = 8'h00;
mem[16'h2403] = 8'h00;
mem[16'h2404] = 8'h42;
mem[16'h2405] = 8'h00;
mem[16'h2406] = 8'h00;
mem[16'h2407] = 8'h00;
mem[16'h2408] = 8'h00;
mem[16'h2409] = 8'h00;
mem[16'h240A] = 8'h42;
mem[16'h240B] = 8'h42;
mem[16'h240C] = 8'h42;
mem[16'h240D] = 8'h42;
mem[16'h240E] = 8'h42;
mem[16'h240F] = 8'h42;
mem[16'h2410] = 8'h00;
mem[16'h2411] = 8'h00;
mem[16'h2412] = 8'h00;
mem[16'h2413] = 8'h00;
mem[16'h2414] = 8'h44;
mem[16'h2415] = 8'h00;
mem[16'h2416] = 8'h00;
mem[16'h2417] = 8'h00;
mem[16'h2418] = 8'h00;
mem[16'h2419] = 8'h42;
mem[16'h241A] = 8'h00;
mem[16'h241B] = 8'h00;
mem[16'h241C] = 8'h00;
mem[16'h241D] = 8'h00;
mem[16'h241E] = 8'h00;
mem[16'h241F] = 8'h42;
mem[16'h2420] = 8'h42;
mem[16'h2421] = 8'h42;
mem[16'h2422] = 8'h42;
mem[16'h2423] = 8'h42;
mem[16'h2424] = 8'h42;
mem[16'h2425] = 8'h00;
mem[16'h2426] = 8'h00;
mem[16'h2427] = 8'h00;
mem[16'h2428] = 8'hD5;
mem[16'h2429] = 8'hAA;
mem[16'h242A] = 8'hD5;
mem[16'h242B] = 8'hAA;
mem[16'h242C] = 8'hD5;
mem[16'h242D] = 8'hD6;
mem[16'h242E] = 8'hAA;
mem[16'h242F] = 8'hD5;
mem[16'h2430] = 8'hAA;
mem[16'h2431] = 8'hD5;
mem[16'h2432] = 8'hAA;
mem[16'h2433] = 8'hB5;
mem[16'h2434] = 8'hD5;
mem[16'h2435] = 8'hAA;
mem[16'h2436] = 8'hD5;
mem[16'h2437] = 8'hAA;
mem[16'h2438] = 8'hD5;
mem[16'h2439] = 8'hDA;
mem[16'h243A] = 8'hAA;
mem[16'h243B] = 8'hD5;
mem[16'h243C] = 8'hAA;
mem[16'h243D] = 8'hD5;
mem[16'h243E] = 8'hAA;
mem[16'h243F] = 8'hD5;
mem[16'h2440] = 8'hD5;
mem[16'h2441] = 8'hAA;
mem[16'h2442] = 8'hD5;
mem[16'h2443] = 8'hAA;
mem[16'h2444] = 8'hB5;
mem[16'h2445] = 8'hD5;
mem[16'h2446] = 8'hAA;
mem[16'h2447] = 8'hD5;
mem[16'h2448] = 8'hAA;
mem[16'h2449] = 8'hD5;
mem[16'h244A] = 8'hAA;
mem[16'h244B] = 8'hAB;
mem[16'h244C] = 8'h85;
mem[16'h244D] = 8'h00;
mem[16'h244E] = 8'h00;
mem[16'h244F] = 8'h00;
mem[16'h2450] = 8'h00;
mem[16'h2451] = 8'hF0;
mem[16'h2452] = 8'hC0;
mem[16'h2453] = 8'h83;
mem[16'h2454] = 8'h00;
mem[16'h2455] = 8'h00;
mem[16'h2456] = 8'h00;
mem[16'h2457] = 8'h00;
mem[16'h2458] = 8'h00;
mem[16'h2459] = 8'h00;
mem[16'h245A] = 8'h00;
mem[16'h245B] = 8'h00;
mem[16'h245C] = 8'h00;
mem[16'h245D] = 8'h00;
mem[16'h245E] = 8'h00;
mem[16'h245F] = 8'h00;
mem[16'h2460] = 8'h00;
mem[16'h2461] = 8'h00;
mem[16'h2462] = 8'h00;
mem[16'h2463] = 8'h00;
mem[16'h2464] = 8'h00;
mem[16'h2465] = 8'h00;
mem[16'h2466] = 8'h00;
mem[16'h2467] = 8'h00;
mem[16'h2468] = 8'h00;
mem[16'h2469] = 8'h00;
mem[16'h246A] = 8'h00;
mem[16'h246B] = 8'h00;
mem[16'h246C] = 8'h00;
mem[16'h246D] = 8'h00;
mem[16'h246E] = 8'h00;
mem[16'h246F] = 8'h00;
mem[16'h2470] = 8'h00;
mem[16'h2471] = 8'h00;
mem[16'h2472] = 8'h00;
mem[16'h2473] = 8'h00;
mem[16'h2474] = 8'h00;
mem[16'h2475] = 8'h00;
mem[16'h2476] = 8'h00;
mem[16'h2477] = 8'h2A;
mem[16'h2478] = 8'h00;
mem[16'h2479] = 8'h00;
mem[16'h247A] = 8'h00;
mem[16'h247B] = 8'h00;
mem[16'h247C] = 8'h00;
mem[16'h247D] = 8'h00;
mem[16'h247E] = 8'h00;
mem[16'h247F] = 8'h00;
mem[16'h2480] = 8'h0A;
mem[16'h2481] = 8'h51;
mem[16'h2482] = 8'h2A;
mem[16'h2483] = 8'hAA;
mem[16'h2484] = 8'hD5;
mem[16'h2485] = 8'h45;
mem[16'h2486] = 8'h2A;
mem[16'h2487] = 8'h51;
mem[16'h2488] = 8'h0A;
mem[16'h2489] = 8'h51;
mem[16'h248A] = 8'hD5;
mem[16'h248B] = 8'hAA;
mem[16'h248C] = 8'h28;
mem[16'h248D] = 8'h45;
mem[16'h248E] = 8'h2A;
mem[16'h248F] = 8'h51;
mem[16'h2490] = 8'hD5;
mem[16'h2491] = 8'hAA;
mem[16'h2492] = 8'h2A;
mem[16'h2493] = 8'h10;
mem[16'h2494] = 8'h28;
mem[16'h2495] = 8'h45;
mem[16'h2496] = 8'h2A;
mem[16'h2497] = 8'hAA;
mem[16'h2498] = 8'hD5;
mem[16'h2499] = 8'h51;
mem[16'h249A] = 8'h2A;
mem[16'h249B] = 8'h10;
mem[16'h249C] = 8'h28;
mem[16'h249D] = 8'hAA;
mem[16'h249E] = 8'hD5;
mem[16'h249F] = 8'h51;
mem[16'h24A0] = 8'h0A;
mem[16'h24A1] = 8'h51;
mem[16'h24A2] = 8'h2A;
mem[16'h24A3] = 8'h10;
mem[16'h24A4] = 8'h08;
mem[16'h24A5] = 8'h00;
mem[16'h24A6] = 8'h74;
mem[16'h24A7] = 8'h17;
mem[16'h24A8] = 8'hD5;
mem[16'h24A9] = 8'hAA;
mem[16'h24AA] = 8'hD5;
mem[16'h24AB] = 8'hAA;
mem[16'h24AC] = 8'hD5;
mem[16'h24AD] = 8'hD6;
mem[16'h24AE] = 8'hAA;
mem[16'h24AF] = 8'hD5;
mem[16'h24B0] = 8'hAA;
mem[16'h24B1] = 8'hD5;
mem[16'h24B2] = 8'hAA;
mem[16'h24B3] = 8'hB5;
mem[16'h24B4] = 8'hD5;
mem[16'h24B5] = 8'hAA;
mem[16'h24B6] = 8'hD5;
mem[16'h24B7] = 8'hAA;
mem[16'h24B8] = 8'hD5;
mem[16'h24B9] = 8'hDA;
mem[16'h24BA] = 8'hAA;
mem[16'h24BB] = 8'hD5;
mem[16'h24BC] = 8'hAA;
mem[16'h24BD] = 8'hD5;
mem[16'h24BE] = 8'hAA;
mem[16'h24BF] = 8'hD5;
mem[16'h24C0] = 8'hD5;
mem[16'h24C1] = 8'hAA;
mem[16'h24C2] = 8'hD5;
mem[16'h24C3] = 8'hAA;
mem[16'h24C4] = 8'hB5;
mem[16'h24C5] = 8'hD5;
mem[16'h24C6] = 8'hAA;
mem[16'h24C7] = 8'hD5;
mem[16'h24C8] = 8'hAA;
mem[16'h24C9] = 8'hD5;
mem[16'h24CA] = 8'hAA;
mem[16'h24CB] = 8'hAB;
mem[16'h24CC] = 8'h85;
mem[16'h24CD] = 8'h00;
mem[16'h24CE] = 8'h00;
mem[16'h24CF] = 8'h2A;
mem[16'h24D0] = 8'h00;
mem[16'h24D1] = 8'h00;
mem[16'h24D2] = 8'h00;
mem[16'h24D3] = 8'h00;
mem[16'h24D4] = 8'h00;
mem[16'h24D5] = 8'h56;
mem[16'h24D6] = 8'h2A;
mem[16'h24D7] = 8'h0F;
mem[16'h24D8] = 8'h00;
mem[16'h24D9] = 8'h00;
mem[16'h24DA] = 8'h00;
mem[16'h24DB] = 8'h00;
mem[16'h24DC] = 8'h00;
mem[16'h24DD] = 8'h00;
mem[16'h24DE] = 8'h00;
mem[16'h24DF] = 8'h00;
mem[16'h24E0] = 8'h00;
mem[16'h24E1] = 8'h56;
mem[16'h24E2] = 8'h2A;
mem[16'h24E3] = 8'h0F;
mem[16'h24E4] = 8'h00;
mem[16'h24E5] = 8'h00;
mem[16'h24E6] = 8'h00;
mem[16'h24E7] = 8'h00;
mem[16'h24E8] = 8'h00;
mem[16'h24E9] = 8'h00;
mem[16'h24EA] = 8'h00;
mem[16'h24EB] = 8'h00;
mem[16'h24EC] = 8'h00;
mem[16'h24ED] = 8'h56;
mem[16'h24EE] = 8'h2A;
mem[16'h24EF] = 8'h0F;
mem[16'h24F0] = 8'h00;
mem[16'h24F1] = 8'h00;
mem[16'h24F2] = 8'h00;
mem[16'h24F3] = 8'h00;
mem[16'h24F4] = 8'h00;
mem[16'h24F5] = 8'h00;
mem[16'h24F6] = 8'h00;
mem[16'h24F7] = 8'h2A;
mem[16'h24F8] = 8'h00;
mem[16'h24F9] = 8'h00;
mem[16'h24FA] = 8'h00;
mem[16'h24FB] = 8'h00;
mem[16'h24FC] = 8'h00;
mem[16'h24FD] = 8'h00;
mem[16'h24FE] = 8'h00;
mem[16'h24FF] = 8'h00;
mem[16'h2500] = 8'h0A;
mem[16'h2501] = 8'h04;
mem[16'h2502] = 8'h2A;
mem[16'h2503] = 8'hAA;
mem[16'h2504] = 8'hD5;
mem[16'h2505] = 8'h54;
mem[16'h2506] = 8'h22;
mem[16'h2507] = 8'h54;
mem[16'h2508] = 8'h0A;
mem[16'h2509] = 8'h04;
mem[16'h250A] = 8'hD5;
mem[16'h250B] = 8'hAA;
mem[16'h250C] = 8'h2A;
mem[16'h250D] = 8'h54;
mem[16'h250E] = 8'h22;
mem[16'h250F] = 8'h54;
mem[16'h2510] = 8'hD5;
mem[16'h2511] = 8'hAA;
mem[16'h2512] = 8'h2A;
mem[16'h2513] = 8'h51;
mem[16'h2514] = 8'h2A;
mem[16'h2515] = 8'h54;
mem[16'h2516] = 8'h22;
mem[16'h2517] = 8'hAA;
mem[16'h2518] = 8'hD5;
mem[16'h2519] = 8'h04;
mem[16'h251A] = 8'h2A;
mem[16'h251B] = 8'h51;
mem[16'h251C] = 8'h2A;
mem[16'h251D] = 8'hAA;
mem[16'h251E] = 8'hD5;
mem[16'h251F] = 8'h54;
mem[16'h2520] = 8'h0A;
mem[16'h2521] = 8'h04;
mem[16'h2522] = 8'h2A;
mem[16'h2523] = 8'h51;
mem[16'h2524] = 8'h0A;
mem[16'h2525] = 8'h00;
mem[16'h2526] = 8'h40;
mem[16'h2527] = 8'h01;
mem[16'h2528] = 8'hD5;
mem[16'h2529] = 8'hAA;
mem[16'h252A] = 8'hD5;
mem[16'h252B] = 8'hAA;
mem[16'h252C] = 8'hD5;
mem[16'h252D] = 8'hCF;
mem[16'h252E] = 8'hAA;
mem[16'h252F] = 8'hFA;
mem[16'h2530] = 8'hA9;
mem[16'h2531] = 8'hA5;
mem[16'h2532] = 8'h9F;
mem[16'h2533] = 8'hD5;
mem[16'h2534] = 8'hD4;
mem[16'h2535] = 8'hAA;
mem[16'h2536] = 8'hD5;
mem[16'h2537] = 8'hAA;
mem[16'h2538] = 8'hD5;
mem[16'h2539] = 8'hAA;
mem[16'h253A] = 8'hD5;
mem[16'h253B] = 8'hEA;
mem[16'h253C] = 8'hA7;
mem[16'h253D] = 8'h95;
mem[16'h253E] = 8'hFD;
mem[16'h253F] = 8'hD4;
mem[16'h2540] = 8'hD2;
mem[16'h2541] = 8'hCF;
mem[16'h2542] = 8'hAA;
mem[16'h2543] = 8'hAA;
mem[16'h2544] = 8'hD5;
mem[16'h2545] = 8'hAA;
mem[16'h2546] = 8'hD5;
mem[16'h2547] = 8'hAA;
mem[16'h2548] = 8'hD5;
mem[16'h2549] = 8'hAA;
mem[16'h254A] = 8'hD5;
mem[16'h254B] = 8'hAA;
mem[16'h254C] = 8'h85;
mem[16'h254D] = 8'h00;
mem[16'h254E] = 8'h00;
mem[16'h254F] = 8'h2A;
mem[16'h2550] = 8'h00;
mem[16'h2551] = 8'h00;
mem[16'h2552] = 8'h00;
mem[16'h2553] = 8'h00;
mem[16'h2554] = 8'h00;
mem[16'h2555] = 8'h00;
mem[16'h2556] = 8'h00;
mem[16'h2557] = 8'h00;
mem[16'h2558] = 8'h00;
mem[16'h2559] = 8'h00;
mem[16'h255A] = 8'h00;
mem[16'h255B] = 8'h00;
mem[16'h255C] = 8'h00;
mem[16'h255D] = 8'h00;
mem[16'h255E] = 8'h00;
mem[16'h255F] = 8'h00;
mem[16'h2560] = 8'h00;
mem[16'h2561] = 8'h00;
mem[16'h2562] = 8'h00;
mem[16'h2563] = 8'h00;
mem[16'h2564] = 8'h00;
mem[16'h2565] = 8'h00;
mem[16'h2566] = 8'h00;
mem[16'h2567] = 8'h00;
mem[16'h2568] = 8'h00;
mem[16'h2569] = 8'h00;
mem[16'h256A] = 8'h00;
mem[16'h256B] = 8'h00;
mem[16'h256C] = 8'h00;
mem[16'h256D] = 8'h00;
mem[16'h256E] = 8'h00;
mem[16'h256F] = 8'h00;
mem[16'h2570] = 8'h00;
mem[16'h2571] = 8'h00;
mem[16'h2572] = 8'h00;
mem[16'h2573] = 8'h00;
mem[16'h2574] = 8'h00;
mem[16'h2575] = 8'h00;
mem[16'h2576] = 8'h00;
mem[16'h2577] = 8'h2A;
mem[16'h2578] = 8'h00;
mem[16'h2579] = 8'h00;
mem[16'h257A] = 8'h00;
mem[16'h257B] = 8'h00;
mem[16'h257C] = 8'h00;
mem[16'h257D] = 8'h00;
mem[16'h257E] = 8'h00;
mem[16'h257F] = 8'h00;
mem[16'h2580] = 8'hD5;
mem[16'h2581] = 8'hAA;
mem[16'h2582] = 8'hD5;
mem[16'h2583] = 8'hAA;
mem[16'h2584] = 8'hD5;
mem[16'h2585] = 8'hAA;
mem[16'h2586] = 8'hAB;
mem[16'h2587] = 8'hD5;
mem[16'h2588] = 8'hAA;
mem[16'h2589] = 8'hD5;
mem[16'h258A] = 8'hAA;
mem[16'h258B] = 8'hD5;
mem[16'h258C] = 8'hAA;
mem[16'h258D] = 8'hD5;
mem[16'h258E] = 8'hAA;
mem[16'h258F] = 8'hD5;
mem[16'h2590] = 8'hD5;
mem[16'h2591] = 8'hAA;
mem[16'h2592] = 8'hAD;
mem[16'h2593] = 8'hD5;
mem[16'h2594] = 8'hAA;
mem[16'h2595] = 8'hD5;
mem[16'h2596] = 8'hAA;
mem[16'h2597] = 8'hD5;
mem[16'h2598] = 8'hAA;
mem[16'h2599] = 8'hD5;
mem[16'h259A] = 8'hAA;
mem[16'h259B] = 8'hD5;
mem[16'h259C] = 8'hD6;
mem[16'h259D] = 8'hAA;
mem[16'h259E] = 8'hD5;
mem[16'h259F] = 8'hAA;
mem[16'h25A0] = 8'hD5;
mem[16'h25A1] = 8'hAA;
mem[16'h25A2] = 8'hD5;
mem[16'h25A3] = 8'hAA;
mem[16'h25A4] = 8'h85;
mem[16'h25A5] = 8'h00;
mem[16'h25A6] = 8'h7C;
mem[16'h25A7] = 8'h1F;
mem[16'h25A8] = 8'hD5;
mem[16'h25A9] = 8'hAA;
mem[16'h25AA] = 8'hD5;
mem[16'h25AB] = 8'hAA;
mem[16'h25AC] = 8'hD5;
mem[16'h25AD] = 8'hAA;
mem[16'h25AE] = 8'hD5;
mem[16'h25AF] = 8'hAA;
mem[16'h25B0] = 8'hD5;
mem[16'h25B1] = 8'hAA;
mem[16'h25B2] = 8'hD5;
mem[16'h25B3] = 8'hAA;
mem[16'h25B4] = 8'hD5;
mem[16'h25B5] = 8'hAA;
mem[16'h25B6] = 8'hD5;
mem[16'h25B7] = 8'hAA;
mem[16'h25B8] = 8'hD5;
mem[16'h25B9] = 8'hAA;
mem[16'h25BA] = 8'hD5;
mem[16'h25BB] = 8'hAA;
mem[16'h25BC] = 8'hD5;
mem[16'h25BD] = 8'hAA;
mem[16'h25BE] = 8'hD5;
mem[16'h25BF] = 8'hAA;
mem[16'h25C0] = 8'hD5;
mem[16'h25C1] = 8'hAA;
mem[16'h25C2] = 8'hD5;
mem[16'h25C3] = 8'hAA;
mem[16'h25C4] = 8'hD5;
mem[16'h25C5] = 8'hAA;
mem[16'h25C6] = 8'hD5;
mem[16'h25C7] = 8'hAA;
mem[16'h25C8] = 8'hD5;
mem[16'h25C9] = 8'hAA;
mem[16'h25CA] = 8'hD5;
mem[16'h25CB] = 8'hAA;
mem[16'h25CC] = 8'h85;
mem[16'h25CD] = 8'h00;
mem[16'h25CE] = 8'h00;
mem[16'h25CF] = 8'h2A;
mem[16'h25D0] = 8'h00;
mem[16'h25D1] = 8'hA8;
mem[16'h25D2] = 8'h95;
mem[16'h25D3] = 8'h81;
mem[16'h25D4] = 8'h00;
mem[16'h25D5] = 8'h00;
mem[16'h25D6] = 8'h00;
mem[16'h25D7] = 8'h00;
mem[16'h25D8] = 8'h00;
mem[16'h25D9] = 8'h00;
mem[16'h25DA] = 8'h00;
mem[16'h25DB] = 8'hC0;
mem[16'h25DC] = 8'hAA;
mem[16'h25DD] = 8'h89;
mem[16'h25DE] = 8'h00;
mem[16'h25DF] = 8'h00;
mem[16'h25E0] = 8'h00;
mem[16'h25E1] = 8'h00;
mem[16'h25E2] = 8'h00;
mem[16'h25E3] = 8'h00;
mem[16'h25E4] = 8'h00;
mem[16'h25E5] = 8'h00;
mem[16'h25E6] = 8'hD4;
mem[16'h25E7] = 8'hCA;
mem[16'h25E8] = 8'h80;
mem[16'h25E9] = 8'h00;
mem[16'h25EA] = 8'h00;
mem[16'h25EB] = 8'h00;
mem[16'h25EC] = 8'h00;
mem[16'h25ED] = 8'h00;
mem[16'h25EE] = 8'h00;
mem[16'h25EF] = 8'h00;
mem[16'h25F0] = 8'h00;
mem[16'h25F1] = 8'h00;
mem[16'h25F2] = 8'h00;
mem[16'h25F3] = 8'h00;
mem[16'h25F4] = 8'h00;
mem[16'h25F5] = 8'h00;
mem[16'h25F6] = 8'h00;
mem[16'h25F7] = 8'h2A;
mem[16'h25F8] = 8'h00;
mem[16'h25F9] = 8'h00;
mem[16'h25FA] = 8'h00;
mem[16'h25FB] = 8'h00;
mem[16'h25FC] = 8'h00;
mem[16'h25FD] = 8'h00;
mem[16'h25FE] = 8'h00;
mem[16'h25FF] = 8'h00;
mem[16'h2600] = 8'hD5;
mem[16'h2601] = 8'hAA;
mem[16'h2602] = 8'hD5;
mem[16'h2603] = 8'hAA;
mem[16'h2604] = 8'hD5;
mem[16'h2605] = 8'hAA;
mem[16'h2606] = 8'hD5;
mem[16'h2607] = 8'hAA;
mem[16'h2608] = 8'hD5;
mem[16'h2609] = 8'hAA;
mem[16'h260A] = 8'hD5;
mem[16'h260B] = 8'hAA;
mem[16'h260C] = 8'hD5;
mem[16'h260D] = 8'hAA;
mem[16'h260E] = 8'hD5;
mem[16'h260F] = 8'hAA;
mem[16'h2610] = 8'hD5;
mem[16'h2611] = 8'hAA;
mem[16'h2612] = 8'hD5;
mem[16'h2613] = 8'hAA;
mem[16'h2614] = 8'hD5;
mem[16'h2615] = 8'hAA;
mem[16'h2616] = 8'hD5;
mem[16'h2617] = 8'hAA;
mem[16'h2618] = 8'hD5;
mem[16'h2619] = 8'hAA;
mem[16'h261A] = 8'hD5;
mem[16'h261B] = 8'hAA;
mem[16'h261C] = 8'hD5;
mem[16'h261D] = 8'hAA;
mem[16'h261E] = 8'hD5;
mem[16'h261F] = 8'hAA;
mem[16'h2620] = 8'hD5;
mem[16'h2621] = 8'hAA;
mem[16'h2622] = 8'hD5;
mem[16'h2623] = 8'hAA;
mem[16'h2624] = 8'h85;
mem[16'h2625] = 8'h00;
mem[16'h2626] = 8'h60;
mem[16'h2627] = 8'h03;
mem[16'h2628] = 8'h02;
mem[16'h2629] = 8'h55;
mem[16'h262A] = 8'h28;
mem[16'h262B] = 8'h15;
mem[16'h262C] = 8'h2A;
mem[16'h262D] = 8'h11;
mem[16'h262E] = 8'h2A;
mem[16'h262F] = 8'h05;
mem[16'h2630] = 8'h02;
mem[16'h2631] = 8'h55;
mem[16'h2632] = 8'h28;
mem[16'h2633] = 8'h15;
mem[16'h2634] = 8'h2A;
mem[16'h2635] = 8'h11;
mem[16'h2636] = 8'h2A;
mem[16'h2637] = 8'h05;
mem[16'h2638] = 8'h02;
mem[16'h2639] = 8'h55;
mem[16'h263A] = 8'h28;
mem[16'h263B] = 8'h15;
mem[16'h263C] = 8'h2A;
mem[16'h263D] = 8'h11;
mem[16'h263E] = 8'h2A;
mem[16'h263F] = 8'h05;
mem[16'h2640] = 8'h02;
mem[16'h2641] = 8'h55;
mem[16'h2642] = 8'h28;
mem[16'h2643] = 8'h15;
mem[16'h2644] = 8'h2A;
mem[16'h2645] = 8'h11;
mem[16'h2646] = 8'h2A;
mem[16'h2647] = 8'h05;
mem[16'h2648] = 8'h02;
mem[16'h2649] = 8'h55;
mem[16'h264A] = 8'h28;
mem[16'h264B] = 8'h15;
mem[16'h264C] = 8'h0A;
mem[16'h264D] = 8'h00;
mem[16'h264E] = 8'h00;
mem[16'h264F] = 8'h2A;
mem[16'h2650] = 8'h00;
mem[16'h2651] = 8'h00;
mem[16'h2652] = 8'h00;
mem[16'h2653] = 8'h00;
mem[16'h2654] = 8'h00;
mem[16'h2655] = 8'h00;
mem[16'h2656] = 8'h00;
mem[16'h2657] = 8'h00;
mem[16'h2658] = 8'h00;
mem[16'h2659] = 8'h00;
mem[16'h265A] = 8'h00;
mem[16'h265B] = 8'h00;
mem[16'h265C] = 8'h00;
mem[16'h265D] = 8'h00;
mem[16'h265E] = 8'h00;
mem[16'h265F] = 8'h00;
mem[16'h2660] = 8'h00;
mem[16'h2661] = 8'h00;
mem[16'h2662] = 8'h00;
mem[16'h2663] = 8'h00;
mem[16'h2664] = 8'h00;
mem[16'h2665] = 8'h00;
mem[16'h2666] = 8'h00;
mem[16'h2667] = 8'h00;
mem[16'h2668] = 8'h00;
mem[16'h2669] = 8'h00;
mem[16'h266A] = 8'h00;
mem[16'h266B] = 8'h00;
mem[16'h266C] = 8'h00;
mem[16'h266D] = 8'h00;
mem[16'h266E] = 8'h00;
mem[16'h266F] = 8'h00;
mem[16'h2670] = 8'h00;
mem[16'h2671] = 8'h00;
mem[16'h2672] = 8'h00;
mem[16'h2673] = 8'h00;
mem[16'h2674] = 8'h00;
mem[16'h2675] = 8'h00;
mem[16'h2676] = 8'h00;
mem[16'h2677] = 8'h2A;
mem[16'h2678] = 8'h00;
mem[16'h2679] = 8'h00;
mem[16'h267A] = 8'h00;
mem[16'h267B] = 8'h00;
mem[16'h267C] = 8'h00;
mem[16'h267D] = 8'h00;
mem[16'h267E] = 8'h00;
mem[16'h267F] = 8'h00;
mem[16'h2680] = 8'hFD;
mem[16'h2681] = 8'hD4;
mem[16'h2682] = 8'hD2;
mem[16'h2683] = 8'hCF;
mem[16'h2684] = 8'hAA;
mem[16'h2685] = 8'hAA;
mem[16'h2686] = 8'hD5;
mem[16'h2687] = 8'hAA;
mem[16'h2688] = 8'hF5;
mem[16'h2689] = 8'hD3;
mem[16'h268A] = 8'hCA;
mem[16'h268B] = 8'hBE;
mem[16'h268C] = 8'hAA;
mem[16'h268D] = 8'hA9;
mem[16'h268E] = 8'hD5;
mem[16'h268F] = 8'hAA;
mem[16'h2690] = 8'hD5;
mem[16'h2691] = 8'hCF;
mem[16'h2692] = 8'hAA;
mem[16'h2693] = 8'hFA;
mem[16'h2694] = 8'hA9;
mem[16'h2695] = 8'hA5;
mem[16'h2696] = 8'hD5;
mem[16'h2697] = 8'hAA;
mem[16'h2698] = 8'hD5;
mem[16'h2699] = 8'hBE;
mem[16'h269A] = 8'hAA;
mem[16'h269B] = 8'hE9;
mem[16'h269C] = 8'hA7;
mem[16'h269D] = 8'h95;
mem[16'h269E] = 8'hD5;
mem[16'h269F] = 8'hAA;
mem[16'h26A0] = 8'hD5;
mem[16'h26A1] = 8'hAA;
mem[16'h26A2] = 8'hD5;
mem[16'h26A3] = 8'hAA;
mem[16'h26A4] = 8'h85;
mem[16'h26A5] = 8'h00;
mem[16'h26A6] = 8'h0E;
mem[16'h26A7] = 8'h38;
mem[16'h26A8] = 8'h00;
mem[16'h26A9] = 8'h00;
mem[16'h26AA] = 8'h00;
mem[16'h26AB] = 8'h00;
mem[16'h26AC] = 8'h00;
mem[16'h26AD] = 8'h00;
mem[16'h26AE] = 8'h00;
mem[16'h26AF] = 8'h00;
mem[16'h26B0] = 8'h00;
mem[16'h26B1] = 8'h00;
mem[16'h26B2] = 8'h00;
mem[16'h26B3] = 8'h00;
mem[16'h26B4] = 8'h00;
mem[16'h26B5] = 8'h00;
mem[16'h26B6] = 8'h00;
mem[16'h26B7] = 8'h00;
mem[16'h26B8] = 8'h00;
mem[16'h26B9] = 8'h00;
mem[16'h26BA] = 8'h00;
mem[16'h26BB] = 8'h00;
mem[16'h26BC] = 8'h00;
mem[16'h26BD] = 8'h00;
mem[16'h26BE] = 8'h00;
mem[16'h26BF] = 8'h00;
mem[16'h26C0] = 8'h00;
mem[16'h26C1] = 8'h00;
mem[16'h26C2] = 8'h00;
mem[16'h26C3] = 8'h00;
mem[16'h26C4] = 8'h00;
mem[16'h26C5] = 8'h00;
mem[16'h26C6] = 8'h00;
mem[16'h26C7] = 8'h00;
mem[16'h26C8] = 8'h00;
mem[16'h26C9] = 8'h00;
mem[16'h26CA] = 8'h00;
mem[16'h26CB] = 8'h00;
mem[16'h26CC] = 8'h00;
mem[16'h26CD] = 8'h00;
mem[16'h26CE] = 8'h00;
mem[16'h26CF] = 8'h2A;
mem[16'h26D0] = 8'h00;
mem[16'h26D1] = 8'h00;
mem[16'h26D2] = 8'h00;
mem[16'h26D3] = 8'h00;
mem[16'h26D4] = 8'h56;
mem[16'h26D5] = 8'h2A;
mem[16'h26D6] = 8'h03;
mem[16'h26D7] = 8'h00;
mem[16'h26D8] = 8'h00;
mem[16'h26D9] = 8'h00;
mem[16'h26DA] = 8'h00;
mem[16'h26DB] = 8'h00;
mem[16'h26DC] = 8'h00;
mem[16'h26DD] = 8'h00;
mem[16'h26DE] = 8'h00;
mem[16'h26DF] = 8'h00;
mem[16'h26E0] = 8'h00;
mem[16'h26E1] = 8'h00;
mem[16'h26E2] = 8'h56;
mem[16'h26E3] = 8'h2A;
mem[16'h26E4] = 8'h03;
mem[16'h26E5] = 8'h00;
mem[16'h26E6] = 8'h00;
mem[16'h26E7] = 8'h00;
mem[16'h26E8] = 8'h00;
mem[16'h26E9] = 8'h00;
mem[16'h26EA] = 8'h00;
mem[16'h26EB] = 8'h00;
mem[16'h26EC] = 8'h00;
mem[16'h26ED] = 8'h00;
mem[16'h26EE] = 8'h00;
mem[16'h26EF] = 8'h00;
mem[16'h26F0] = 8'h56;
mem[16'h26F1] = 8'h2A;
mem[16'h26F2] = 8'h03;
mem[16'h26F3] = 8'h00;
mem[16'h26F4] = 8'h00;
mem[16'h26F5] = 8'h00;
mem[16'h26F6] = 8'h00;
mem[16'h26F7] = 8'h2A;
mem[16'h26F8] = 8'h00;
mem[16'h26F9] = 8'h00;
mem[16'h26FA] = 8'h00;
mem[16'h26FB] = 8'h00;
mem[16'h26FC] = 8'h00;
mem[16'h26FD] = 8'h00;
mem[16'h26FE] = 8'h00;
mem[16'h26FF] = 8'h00;
mem[16'h2700] = 8'hD5;
mem[16'h2701] = 8'hAA;
mem[16'h2702] = 8'hD5;
mem[16'h2703] = 8'hAA;
mem[16'h2704] = 8'hD5;
mem[16'h2705] = 8'hAA;
mem[16'h2706] = 8'hD5;
mem[16'h2707] = 8'hAA;
mem[16'h2708] = 8'hD5;
mem[16'h2709] = 8'hAA;
mem[16'h270A] = 8'hD5;
mem[16'h270B] = 8'hAA;
mem[16'h270C] = 8'hD5;
mem[16'h270D] = 8'hAA;
mem[16'h270E] = 8'hD5;
mem[16'h270F] = 8'hAA;
mem[16'h2710] = 8'hD5;
mem[16'h2711] = 8'hAA;
mem[16'h2712] = 8'hD5;
mem[16'h2713] = 8'hAA;
mem[16'h2714] = 8'hD5;
mem[16'h2715] = 8'hAA;
mem[16'h2716] = 8'hD5;
mem[16'h2717] = 8'hAA;
mem[16'h2718] = 8'hD5;
mem[16'h2719] = 8'hAA;
mem[16'h271A] = 8'hD5;
mem[16'h271B] = 8'hAA;
mem[16'h271C] = 8'hD5;
mem[16'h271D] = 8'hAA;
mem[16'h271E] = 8'hD5;
mem[16'h271F] = 8'hAA;
mem[16'h2720] = 8'hD5;
mem[16'h2721] = 8'hAA;
mem[16'h2722] = 8'hD5;
mem[16'h2723] = 8'hAA;
mem[16'h2724] = 8'h85;
mem[16'h2725] = 8'h00;
mem[16'h2726] = 8'h60;
mem[16'h2727] = 8'h03;
mem[16'h2728] = 8'h00;
mem[16'h2729] = 8'h00;
mem[16'h272A] = 8'h1D;
mem[16'h272B] = 8'h55;
mem[16'h272C] = 8'h0A;
mem[16'h272D] = 8'h00;
mem[16'h272E] = 8'h00;
mem[16'h272F] = 8'h00;
mem[16'h2730] = 8'h00;
mem[16'h2731] = 8'h00;
mem[16'h2732] = 8'h00;
mem[16'h2733] = 8'h00;
mem[16'h2734] = 8'h00;
mem[16'h2735] = 8'h00;
mem[16'h2736] = 8'h00;
mem[16'h2737] = 8'h00;
mem[16'h2738] = 8'h1D;
mem[16'h2739] = 8'h55;
mem[16'h273A] = 8'h0A;
mem[16'h273B] = 8'h00;
mem[16'h273C] = 8'h00;
mem[16'h273D] = 8'h00;
mem[16'h273E] = 8'h00;
mem[16'h273F] = 8'h00;
mem[16'h2740] = 8'h00;
mem[16'h2741] = 8'h00;
mem[16'h2742] = 8'h00;
mem[16'h2743] = 8'h00;
mem[16'h2744] = 8'h00;
mem[16'h2745] = 8'h00;
mem[16'h2746] = 8'h00;
mem[16'h2747] = 8'h00;
mem[16'h2748] = 8'h00;
mem[16'h2749] = 8'h00;
mem[16'h274A] = 8'h00;
mem[16'h274B] = 8'h00;
mem[16'h274C] = 8'h00;
mem[16'h274D] = 8'h00;
mem[16'h274E] = 8'h00;
mem[16'h274F] = 8'h2A;
mem[16'h2750] = 8'h28;
mem[16'h2751] = 8'h15;
mem[16'h2752] = 8'h08;
mem[16'h2753] = 8'h54;
mem[16'h2754] = 8'h22;
mem[16'h2755] = 8'h55;
mem[16'h2756] = 8'h28;
mem[16'h2757] = 8'h45;
mem[16'h2758] = 8'h28;
mem[16'h2759] = 8'h15;
mem[16'h275A] = 8'h08;
mem[16'h275B] = 8'h54;
mem[16'h275C] = 8'h22;
mem[16'h275D] = 8'h55;
mem[16'h275E] = 8'h28;
mem[16'h275F] = 8'h45;
mem[16'h2760] = 8'h28;
mem[16'h2761] = 8'h15;
mem[16'h2762] = 8'h60;
mem[16'h2763] = 8'h03;
mem[16'h2764] = 8'h22;
mem[16'h2765] = 8'h55;
mem[16'h2766] = 8'h28;
mem[16'h2767] = 8'h45;
mem[16'h2768] = 8'h28;
mem[16'h2769] = 8'h15;
mem[16'h276A] = 8'h08;
mem[16'h276B] = 8'h54;
mem[16'h276C] = 8'h22;
mem[16'h276D] = 8'h55;
mem[16'h276E] = 8'h28;
mem[16'h276F] = 8'h45;
mem[16'h2770] = 8'h28;
mem[16'h2771] = 8'h15;
mem[16'h2772] = 8'h08;
mem[16'h2773] = 8'h54;
mem[16'h2774] = 8'h02;
mem[16'h2775] = 8'h00;
mem[16'h2776] = 8'h00;
mem[16'h2777] = 8'h2A;
mem[16'h2778] = 8'h00;
mem[16'h2779] = 8'h00;
mem[16'h277A] = 8'h00;
mem[16'h277B] = 8'h00;
mem[16'h277C] = 8'h00;
mem[16'h277D] = 8'h00;
mem[16'h277E] = 8'h00;
mem[16'h277F] = 8'h00;
mem[16'h2780] = 8'hAB;
mem[16'h2781] = 8'hAD;
mem[16'h2782] = 8'hD5;
mem[16'h2783] = 8'hAA;
mem[16'h2784] = 8'hD5;
mem[16'h2785] = 8'hAA;
mem[16'h2786] = 8'hD5;
mem[16'h2787] = 8'hAA;
mem[16'h2788] = 8'hD5;
mem[16'h2789] = 8'hAA;
mem[16'h278A] = 8'hD5;
mem[16'h278B] = 8'hD5;
mem[16'h278C] = 8'hAA;
mem[16'h278D] = 8'hD5;
mem[16'h278E] = 8'hAA;
mem[16'h278F] = 8'hD5;
mem[16'h2790] = 8'hAA;
mem[16'h2791] = 8'hD5;
mem[16'h2792] = 8'hAA;
mem[16'h2793] = 8'hD5;
mem[16'h2794] = 8'hAA;
mem[16'h2795] = 8'hD5;
mem[16'h2796] = 8'hAA;
mem[16'h2797] = 8'hD5;
mem[16'h2798] = 8'hAA;
mem[16'h2799] = 8'hD5;
mem[16'h279A] = 8'hD5;
mem[16'h279B] = 8'hAA;
mem[16'h279C] = 8'hD5;
mem[16'h279D] = 8'hAA;
mem[16'h279E] = 8'hD5;
mem[16'h279F] = 8'hAA;
mem[16'h27A0] = 8'hD5;
mem[16'h27A1] = 8'hAA;
mem[16'h27A2] = 8'hD5;
mem[16'h27A3] = 8'hAA;
mem[16'h27A4] = 8'h85;
mem[16'h27A5] = 8'h00;
mem[16'h27A6] = 8'h00;
mem[16'h27A7] = 8'h00;
mem[16'h27A8] = 8'h00;
mem[16'h27A9] = 8'h00;
mem[16'h27AA] = 8'h00;
mem[16'h27AB] = 8'h00;
mem[16'h27AC] = 8'h00;
mem[16'h27AD] = 8'h00;
mem[16'h27AE] = 8'h00;
mem[16'h27AF] = 8'h00;
mem[16'h27B0] = 8'h00;
mem[16'h27B1] = 8'h00;
mem[16'h27B2] = 8'h00;
mem[16'h27B3] = 8'h00;
mem[16'h27B4] = 8'h00;
mem[16'h27B5] = 8'h00;
mem[16'h27B6] = 8'h00;
mem[16'h27B7] = 8'h00;
mem[16'h27B8] = 8'h00;
mem[16'h27B9] = 8'h00;
mem[16'h27BA] = 8'h00;
mem[16'h27BB] = 8'h00;
mem[16'h27BC] = 8'h00;
mem[16'h27BD] = 8'h00;
mem[16'h27BE] = 8'h00;
mem[16'h27BF] = 8'h00;
mem[16'h27C0] = 8'h00;
mem[16'h27C1] = 8'h00;
mem[16'h27C2] = 8'h00;
mem[16'h27C3] = 8'h00;
mem[16'h27C4] = 8'h00;
mem[16'h27C5] = 8'h00;
mem[16'h27C6] = 8'h00;
mem[16'h27C7] = 8'h00;
mem[16'h27C8] = 8'h00;
mem[16'h27C9] = 8'h00;
mem[16'h27CA] = 8'h00;
mem[16'h27CB] = 8'h00;
mem[16'h27CC] = 8'h00;
mem[16'h27CD] = 8'h00;
mem[16'h27CE] = 8'h00;
mem[16'h27CF] = 8'h2A;
mem[16'h27D0] = 8'h28;
mem[16'h27D1] = 8'h15;
mem[16'h27D2] = 8'h08;
mem[16'h27D3] = 8'h54;
mem[16'h27D4] = 8'h22;
mem[16'h27D5] = 8'h55;
mem[16'h27D6] = 8'h28;
mem[16'h27D7] = 8'h45;
mem[16'h27D8] = 8'h28;
mem[16'h27D9] = 8'h15;
mem[16'h27DA] = 8'h08;
mem[16'h27DB] = 8'h54;
mem[16'h27DC] = 8'h22;
mem[16'h27DD] = 8'h55;
mem[16'h27DE] = 8'h28;
mem[16'h27DF] = 8'h45;
mem[16'h27E0] = 8'h28;
mem[16'h27E1] = 8'h15;
mem[16'h27E2] = 8'h44;
mem[16'h27E3] = 8'h12;
mem[16'h27E4] = 8'h22;
mem[16'h27E5] = 8'h55;
mem[16'h27E6] = 8'h28;
mem[16'h27E7] = 8'h45;
mem[16'h27E8] = 8'h28;
mem[16'h27E9] = 8'h15;
mem[16'h27EA] = 8'h08;
mem[16'h27EB] = 8'h54;
mem[16'h27EC] = 8'h22;
mem[16'h27ED] = 8'h55;
mem[16'h27EE] = 8'h28;
mem[16'h27EF] = 8'h45;
mem[16'h27F0] = 8'h28;
mem[16'h27F1] = 8'h15;
mem[16'h27F2] = 8'h08;
mem[16'h27F3] = 8'h54;
mem[16'h27F4] = 8'h02;
mem[16'h27F5] = 8'h46;
mem[16'h27F6] = 8'h00;
mem[16'h27F7] = 8'h2A;
mem[16'h27F8] = 8'h00;
mem[16'h27F9] = 8'h00;
mem[16'h27FA] = 8'h00;
mem[16'h27FB] = 8'h00;
mem[16'h27FC] = 8'h00;
mem[16'h27FD] = 8'h00;
mem[16'h27FE] = 8'h00;
mem[16'h27FF] = 8'h00;
mem[16'h2800] = 8'h00;
mem[16'h2801] = 8'h42;
mem[16'h2802] = 8'h18;
mem[16'h2803] = 8'h00;
mem[16'h2804] = 8'h02;
mem[16'h2805] = 8'h3C;
mem[16'h2806] = 8'h38;
mem[16'h2807] = 8'h3A;
mem[16'h2808] = 8'h3C;
mem[16'h2809] = 8'h00;
mem[16'h280A] = 8'h42;
mem[16'h280B] = 8'h42;
mem[16'h280C] = 8'h42;
mem[16'h280D] = 8'h42;
mem[16'h280E] = 8'h42;
mem[16'h280F] = 8'h42;
mem[16'h2810] = 8'h00;
mem[16'h2811] = 8'h00;
mem[16'h2812] = 8'h00;
mem[16'h2813] = 8'h00;
mem[16'h2814] = 8'h44;
mem[16'h2815] = 8'h38;
mem[16'h2816] = 8'h42;
mem[16'h2817] = 8'h3A;
mem[16'h2818] = 8'h00;
mem[16'h2819] = 8'h02;
mem[16'h281A] = 8'h3C;
mem[16'h281B] = 8'h38;
mem[16'h281C] = 8'h3A;
mem[16'h281D] = 8'h3C;
mem[16'h281E] = 8'h00;
mem[16'h281F] = 8'h42;
mem[16'h2820] = 8'h42;
mem[16'h2821] = 8'h42;
mem[16'h2822] = 8'h42;
mem[16'h2823] = 8'h42;
mem[16'h2824] = 8'h42;
mem[16'h2825] = 8'h00;
mem[16'h2826] = 8'h00;
mem[16'h2827] = 8'h00;
mem[16'h2828] = 8'hD5;
mem[16'h2829] = 8'hAA;
mem[16'h282A] = 8'hD5;
mem[16'h282B] = 8'hAA;
mem[16'h282C] = 8'hD5;
mem[16'h282D] = 8'hD5;
mem[16'h282E] = 8'hAA;
mem[16'h282F] = 8'hD5;
mem[16'h2830] = 8'hAA;
mem[16'h2831] = 8'hD5;
mem[16'h2832] = 8'hAA;
mem[16'h2833] = 8'hD5;
mem[16'h2834] = 8'hD5;
mem[16'h2835] = 8'hAA;
mem[16'h2836] = 8'hD5;
mem[16'h2837] = 8'hAA;
mem[16'h2838] = 8'hD5;
mem[16'h2839] = 8'hD6;
mem[16'h283A] = 8'hAA;
mem[16'h283B] = 8'hD5;
mem[16'h283C] = 8'hAA;
mem[16'h283D] = 8'hD5;
mem[16'h283E] = 8'hAA;
mem[16'h283F] = 8'hD5;
mem[16'h2840] = 8'hD6;
mem[16'h2841] = 8'hAA;
mem[16'h2842] = 8'hD5;
mem[16'h2843] = 8'hAA;
mem[16'h2844] = 8'hAD;
mem[16'h2845] = 8'hD5;
mem[16'h2846] = 8'hAA;
mem[16'h2847] = 8'hD5;
mem[16'h2848] = 8'hAA;
mem[16'h2849] = 8'hD5;
mem[16'h284A] = 8'hAA;
mem[16'h284B] = 8'hAD;
mem[16'h284C] = 8'h85;
mem[16'h284D] = 8'h00;
mem[16'h284E] = 8'h00;
mem[16'h284F] = 8'h00;
mem[16'h2850] = 8'h00;
mem[16'h2851] = 8'h00;
mem[16'h2852] = 8'h00;
mem[16'h2853] = 8'h00;
mem[16'h2854] = 8'h00;
mem[16'h2855] = 8'h00;
mem[16'h2856] = 8'h00;
mem[16'h2857] = 8'h00;
mem[16'h2858] = 8'h00;
mem[16'h2859] = 8'h00;
mem[16'h285A] = 8'h00;
mem[16'h285B] = 8'h00;
mem[16'h285C] = 8'h00;
mem[16'h285D] = 8'h00;
mem[16'h285E] = 8'h00;
mem[16'h285F] = 8'h00;
mem[16'h2860] = 8'h00;
mem[16'h2861] = 8'h00;
mem[16'h2862] = 8'h00;
mem[16'h2863] = 8'h00;
mem[16'h2864] = 8'h00;
mem[16'h2865] = 8'h00;
mem[16'h2866] = 8'h00;
mem[16'h2867] = 8'h00;
mem[16'h2868] = 8'h00;
mem[16'h2869] = 8'h00;
mem[16'h286A] = 8'h00;
mem[16'h286B] = 8'h00;
mem[16'h286C] = 8'h00;
mem[16'h286D] = 8'h00;
mem[16'h286E] = 8'h00;
mem[16'h286F] = 8'h00;
mem[16'h2870] = 8'h00;
mem[16'h2871] = 8'h00;
mem[16'h2872] = 8'h00;
mem[16'h2873] = 8'h00;
mem[16'h2874] = 8'h00;
mem[16'h2875] = 8'h00;
mem[16'h2876] = 8'h00;
mem[16'h2877] = 8'h2A;
mem[16'h2878] = 8'h00;
mem[16'h2879] = 8'h00;
mem[16'h287A] = 8'h00;
mem[16'h287B] = 8'h00;
mem[16'h287C] = 8'h00;
mem[16'h287D] = 8'h00;
mem[16'h287E] = 8'h00;
mem[16'h287F] = 8'h00;
mem[16'h2880] = 8'h2A;
mem[16'h2881] = 8'h54;
mem[16'h2882] = 8'h0A;
mem[16'h2883] = 8'hAA;
mem[16'h2884] = 8'hD5;
mem[16'h2885] = 8'h55;
mem[16'h2886] = 8'h02;
mem[16'h2887] = 8'h41;
mem[16'h2888] = 8'h2A;
mem[16'h2889] = 8'h54;
mem[16'h288A] = 8'hD5;
mem[16'h288B] = 8'hAA;
mem[16'h288C] = 8'h08;
mem[16'h288D] = 8'h55;
mem[16'h288E] = 8'h02;
mem[16'h288F] = 8'h41;
mem[16'h2890] = 8'hD5;
mem[16'h2891] = 8'hAA;
mem[16'h2892] = 8'h0A;
mem[16'h2893] = 8'h55;
mem[16'h2894] = 8'h08;
mem[16'h2895] = 8'h55;
mem[16'h2896] = 8'h02;
mem[16'h2897] = 8'hAA;
mem[16'h2898] = 8'hD5;
mem[16'h2899] = 8'h54;
mem[16'h289A] = 8'h0A;
mem[16'h289B] = 8'h55;
mem[16'h289C] = 8'h08;
mem[16'h289D] = 8'hAA;
mem[16'h289E] = 8'hD5;
mem[16'h289F] = 8'h41;
mem[16'h28A0] = 8'h2A;
mem[16'h28A1] = 8'h54;
mem[16'h28A2] = 8'h0A;
mem[16'h28A3] = 8'h55;
mem[16'h28A4] = 8'h08;
mem[16'h28A5] = 8'h00;
mem[16'h28A6] = 8'h7C;
mem[16'h28A7] = 8'h1F;
mem[16'h28A8] = 8'hD5;
mem[16'h28A9] = 8'hAA;
mem[16'h28AA] = 8'hD5;
mem[16'h28AB] = 8'hAA;
mem[16'h28AC] = 8'hD5;
mem[16'h28AD] = 8'hAA;
mem[16'h28AE] = 8'hD5;
mem[16'h28AF] = 8'hAA;
mem[16'h28B0] = 8'hD5;
mem[16'h28B1] = 8'hAA;
mem[16'h28B2] = 8'hD5;
mem[16'h28B3] = 8'hAA;
mem[16'h28B4] = 8'hD5;
mem[16'h28B5] = 8'hAA;
mem[16'h28B6] = 8'hD5;
mem[16'h28B7] = 8'hAA;
mem[16'h28B8] = 8'hD5;
mem[16'h28B9] = 8'hAA;
mem[16'h28BA] = 8'hD5;
mem[16'h28BB] = 8'hAA;
mem[16'h28BC] = 8'hD5;
mem[16'h28BD] = 8'hAA;
mem[16'h28BE] = 8'hD5;
mem[16'h28BF] = 8'hAA;
mem[16'h28C0] = 8'hD5;
mem[16'h28C1] = 8'hAA;
mem[16'h28C2] = 8'hD5;
mem[16'h28C3] = 8'hAA;
mem[16'h28C4] = 8'hD5;
mem[16'h28C5] = 8'hAA;
mem[16'h28C6] = 8'hD5;
mem[16'h28C7] = 8'hAA;
mem[16'h28C8] = 8'hD5;
mem[16'h28C9] = 8'hAA;
mem[16'h28CA] = 8'hD5;
mem[16'h28CB] = 8'hAA;
mem[16'h28CC] = 8'h85;
mem[16'h28CD] = 8'h00;
mem[16'h28CE] = 8'h00;
mem[16'h28CF] = 8'h2A;
mem[16'h28D0] = 8'h00;
mem[16'h28D1] = 8'h00;
mem[16'h28D2] = 8'h00;
mem[16'h28D3] = 8'h00;
mem[16'h28D4] = 8'h00;
mem[16'h28D5] = 8'h55;
mem[16'h28D6] = 8'h28;
mem[16'h28D7] = 8'h03;
mem[16'h28D8] = 8'h00;
mem[16'h28D9] = 8'h00;
mem[16'h28DA] = 8'h00;
mem[16'h28DB] = 8'h00;
mem[16'h28DC] = 8'h00;
mem[16'h28DD] = 8'h00;
mem[16'h28DE] = 8'h00;
mem[16'h28DF] = 8'h00;
mem[16'h28E0] = 8'h00;
mem[16'h28E1] = 8'h55;
mem[16'h28E2] = 8'h28;
mem[16'h28E3] = 8'h03;
mem[16'h28E4] = 8'h00;
mem[16'h28E5] = 8'h00;
mem[16'h28E6] = 8'h00;
mem[16'h28E7] = 8'h00;
mem[16'h28E8] = 8'h00;
mem[16'h28E9] = 8'h00;
mem[16'h28EA] = 8'h00;
mem[16'h28EB] = 8'h00;
mem[16'h28EC] = 8'h00;
mem[16'h28ED] = 8'h55;
mem[16'h28EE] = 8'h28;
mem[16'h28EF] = 8'h03;
mem[16'h28F0] = 8'h00;
mem[16'h28F1] = 8'h00;
mem[16'h28F2] = 8'h00;
mem[16'h28F3] = 8'h00;
mem[16'h28F4] = 8'h00;
mem[16'h28F5] = 8'h00;
mem[16'h28F6] = 8'h00;
mem[16'h28F7] = 8'h2A;
mem[16'h28F8] = 8'h00;
mem[16'h28F9] = 8'h00;
mem[16'h28FA] = 8'h00;
mem[16'h28FB] = 8'h00;
mem[16'h28FC] = 8'h00;
mem[16'h28FD] = 8'h00;
mem[16'h28FE] = 8'h00;
mem[16'h28FF] = 8'h00;
mem[16'h2900] = 8'h2A;
mem[16'h2901] = 8'h54;
mem[16'h2902] = 8'h0A;
mem[16'h2903] = 8'hAA;
mem[16'h2904] = 8'hD5;
mem[16'h2905] = 8'h55;
mem[16'h2906] = 8'h02;
mem[16'h2907] = 8'h41;
mem[16'h2908] = 8'h2A;
mem[16'h2909] = 8'h54;
mem[16'h290A] = 8'hD5;
mem[16'h290B] = 8'hAA;
mem[16'h290C] = 8'h08;
mem[16'h290D] = 8'h55;
mem[16'h290E] = 8'h02;
mem[16'h290F] = 8'h41;
mem[16'h2910] = 8'hD5;
mem[16'h2911] = 8'hAA;
mem[16'h2912] = 8'h0A;
mem[16'h2913] = 8'h55;
mem[16'h2914] = 8'h08;
mem[16'h2915] = 8'h55;
mem[16'h2916] = 8'h02;
mem[16'h2917] = 8'hAA;
mem[16'h2918] = 8'hD5;
mem[16'h2919] = 8'h54;
mem[16'h291A] = 8'h0A;
mem[16'h291B] = 8'h55;
mem[16'h291C] = 8'h08;
mem[16'h291D] = 8'hAA;
mem[16'h291E] = 8'hD5;
mem[16'h291F] = 8'h41;
mem[16'h2920] = 8'h2A;
mem[16'h2921] = 8'h54;
mem[16'h2922] = 8'h0A;
mem[16'h2923] = 8'h55;
mem[16'h2924] = 8'h08;
mem[16'h2925] = 8'h00;
mem[16'h2926] = 8'h60;
mem[16'h2927] = 8'h03;
mem[16'h2928] = 8'hD5;
mem[16'h2929] = 8'hAA;
mem[16'h292A] = 8'hD5;
mem[16'h292B] = 8'hAA;
mem[16'h292C] = 8'hD5;
mem[16'h292D] = 8'hCF;
mem[16'h292E] = 8'hAA;
mem[16'h292F] = 8'hFA;
mem[16'h2930] = 8'hA9;
mem[16'h2931] = 8'hA5;
mem[16'h2932] = 8'h9F;
mem[16'h2933] = 8'hD5;
mem[16'h2934] = 8'hD4;
mem[16'h2935] = 8'hAA;
mem[16'h2936] = 8'hD5;
mem[16'h2937] = 8'hAA;
mem[16'h2938] = 8'hD5;
mem[16'h2939] = 8'hAA;
mem[16'h293A] = 8'hD5;
mem[16'h293B] = 8'hEA;
mem[16'h293C] = 8'hA7;
mem[16'h293D] = 8'h95;
mem[16'h293E] = 8'hFD;
mem[16'h293F] = 8'hD4;
mem[16'h2940] = 8'hD2;
mem[16'h2941] = 8'hCF;
mem[16'h2942] = 8'hAA;
mem[16'h2943] = 8'hAA;
mem[16'h2944] = 8'hD5;
mem[16'h2945] = 8'hAA;
mem[16'h2946] = 8'hD5;
mem[16'h2947] = 8'hAA;
mem[16'h2948] = 8'hD5;
mem[16'h2949] = 8'hAA;
mem[16'h294A] = 8'hD5;
mem[16'h294B] = 8'hAA;
mem[16'h294C] = 8'h85;
mem[16'h294D] = 8'h00;
mem[16'h294E] = 8'h00;
mem[16'h294F] = 8'h2A;
mem[16'h2950] = 8'h00;
mem[16'h2951] = 8'h00;
mem[16'h2952] = 8'h00;
mem[16'h2953] = 8'h00;
mem[16'h2954] = 8'h00;
mem[16'h2955] = 8'h00;
mem[16'h2956] = 8'h00;
mem[16'h2957] = 8'h00;
mem[16'h2958] = 8'h00;
mem[16'h2959] = 8'h00;
mem[16'h295A] = 8'h00;
mem[16'h295B] = 8'h00;
mem[16'h295C] = 8'h00;
mem[16'h295D] = 8'h00;
mem[16'h295E] = 8'h00;
mem[16'h295F] = 8'h00;
mem[16'h2960] = 8'h00;
mem[16'h2961] = 8'h00;
mem[16'h2962] = 8'h00;
mem[16'h2963] = 8'h00;
mem[16'h2964] = 8'h00;
mem[16'h2965] = 8'h00;
mem[16'h2966] = 8'h00;
mem[16'h2967] = 8'h00;
mem[16'h2968] = 8'h00;
mem[16'h2969] = 8'h00;
mem[16'h296A] = 8'h00;
mem[16'h296B] = 8'h00;
mem[16'h296C] = 8'h00;
mem[16'h296D] = 8'h00;
mem[16'h296E] = 8'h00;
mem[16'h296F] = 8'h00;
mem[16'h2970] = 8'h00;
mem[16'h2971] = 8'h00;
mem[16'h2972] = 8'h00;
mem[16'h2973] = 8'h00;
mem[16'h2974] = 8'h00;
mem[16'h2975] = 8'h00;
mem[16'h2976] = 8'h00;
mem[16'h2977] = 8'h2A;
mem[16'h2978] = 8'h00;
mem[16'h2979] = 8'h00;
mem[16'h297A] = 8'h00;
mem[16'h297B] = 8'h00;
mem[16'h297C] = 8'h00;
mem[16'h297D] = 8'h00;
mem[16'h297E] = 8'h00;
mem[16'h297F] = 8'h00;
mem[16'h2980] = 8'hD5;
mem[16'h2981] = 8'hAA;
mem[16'h2982] = 8'hD5;
mem[16'h2983] = 8'hAA;
mem[16'h2984] = 8'hD5;
mem[16'h2985] = 8'hAA;
mem[16'h2986] = 8'hAB;
mem[16'h2987] = 8'hD5;
mem[16'h2988] = 8'hAA;
mem[16'h2989] = 8'hD5;
mem[16'h298A] = 8'hAA;
mem[16'h298B] = 8'hD5;
mem[16'h298C] = 8'hAA;
mem[16'h298D] = 8'hD5;
mem[16'h298E] = 8'hAA;
mem[16'h298F] = 8'hD5;
mem[16'h2990] = 8'hD5;
mem[16'h2991] = 8'hAA;
mem[16'h2992] = 8'hAD;
mem[16'h2993] = 8'hD5;
mem[16'h2994] = 8'hAA;
mem[16'h2995] = 8'hD5;
mem[16'h2996] = 8'hAA;
mem[16'h2997] = 8'hD5;
mem[16'h2998] = 8'hAA;
mem[16'h2999] = 8'hD5;
mem[16'h299A] = 8'hAA;
mem[16'h299B] = 8'hD5;
mem[16'h299C] = 8'hD6;
mem[16'h299D] = 8'hAA;
mem[16'h299E] = 8'hD5;
mem[16'h299F] = 8'hAA;
mem[16'h29A0] = 8'hD5;
mem[16'h29A1] = 8'hAA;
mem[16'h29A2] = 8'hD5;
mem[16'h29A3] = 8'hAA;
mem[16'h29A4] = 8'h85;
mem[16'h29A5] = 8'h00;
mem[16'h29A6] = 8'h44;
mem[16'h29A7] = 8'h12;
mem[16'h29A8] = 8'h2A;
mem[16'h29A9] = 8'h45;
mem[16'h29AA] = 8'h2A;
mem[16'h29AB] = 8'h44;
mem[16'h29AC] = 8'h2A;
mem[16'h29AD] = 8'h41;
mem[16'h29AE] = 8'h20;
mem[16'h29AF] = 8'h15;
mem[16'h29B0] = 8'h2A;
mem[16'h29B1] = 8'h45;
mem[16'h29B2] = 8'h2A;
mem[16'h29B3] = 8'h44;
mem[16'h29B4] = 8'h2A;
mem[16'h29B5] = 8'h41;
mem[16'h29B6] = 8'h20;
mem[16'h29B7] = 8'h15;
mem[16'h29B8] = 8'h2A;
mem[16'h29B9] = 8'h45;
mem[16'h29BA] = 8'h2A;
mem[16'h29BB] = 8'h44;
mem[16'h29BC] = 8'h2A;
mem[16'h29BD] = 8'h41;
mem[16'h29BE] = 8'h20;
mem[16'h29BF] = 8'h15;
mem[16'h29C0] = 8'h2A;
mem[16'h29C1] = 8'h45;
mem[16'h29C2] = 8'h2A;
mem[16'h29C3] = 8'h44;
mem[16'h29C4] = 8'h2A;
mem[16'h29C5] = 8'h41;
mem[16'h29C6] = 8'h20;
mem[16'h29C7] = 8'h15;
mem[16'h29C8] = 8'h2A;
mem[16'h29C9] = 8'h45;
mem[16'h29CA] = 8'h2A;
mem[16'h29CB] = 8'h44;
mem[16'h29CC] = 8'h0A;
mem[16'h29CD] = 8'h00;
mem[16'h29CE] = 8'h00;
mem[16'h29CF] = 8'h2A;
mem[16'h29D0] = 8'h00;
mem[16'h29D1] = 8'hA8;
mem[16'h29D2] = 8'hF5;
mem[16'h29D3] = 8'h81;
mem[16'h29D4] = 8'h00;
mem[16'h29D5] = 8'h00;
mem[16'h29D6] = 8'h00;
mem[16'h29D7] = 8'h00;
mem[16'h29D8] = 8'h00;
mem[16'h29D9] = 8'h00;
mem[16'h29DA] = 8'h00;
mem[16'h29DB] = 8'hC0;
mem[16'h29DC] = 8'hAA;
mem[16'h29DD] = 8'h8F;
mem[16'h29DE] = 8'h00;
mem[16'h29DF] = 8'h00;
mem[16'h29E0] = 8'h00;
mem[16'h29E1] = 8'h00;
mem[16'h29E2] = 8'h00;
mem[16'h29E3] = 8'h00;
mem[16'h29E4] = 8'h00;
mem[16'h29E5] = 8'h00;
mem[16'h29E6] = 8'hD4;
mem[16'h29E7] = 8'hFA;
mem[16'h29E8] = 8'h80;
mem[16'h29E9] = 8'h00;
mem[16'h29EA] = 8'h00;
mem[16'h29EB] = 8'h00;
mem[16'h29EC] = 8'h00;
mem[16'h29ED] = 8'h00;
mem[16'h29EE] = 8'h00;
mem[16'h29EF] = 8'h00;
mem[16'h29F0] = 8'h00;
mem[16'h29F1] = 8'h00;
mem[16'h29F2] = 8'h00;
mem[16'h29F3] = 8'h00;
mem[16'h29F4] = 8'h00;
mem[16'h29F5] = 8'h00;
mem[16'h29F6] = 8'h00;
mem[16'h29F7] = 8'h2A;
mem[16'h29F8] = 8'h00;
mem[16'h29F9] = 8'h00;
mem[16'h29FA] = 8'h00;
mem[16'h29FB] = 8'h00;
mem[16'h29FC] = 8'h00;
mem[16'h29FD] = 8'h00;
mem[16'h29FE] = 8'h00;
mem[16'h29FF] = 8'h00;
mem[16'h2A00] = 8'hD5;
mem[16'h2A01] = 8'hAA;
mem[16'h2A02] = 8'hD5;
mem[16'h2A03] = 8'hAA;
mem[16'h2A04] = 8'hD5;
mem[16'h2A05] = 8'hAA;
mem[16'h2A06] = 8'hD5;
mem[16'h2A07] = 8'hAA;
mem[16'h2A08] = 8'hD5;
mem[16'h2A09] = 8'hAA;
mem[16'h2A0A] = 8'hD5;
mem[16'h2A0B] = 8'hAA;
mem[16'h2A0C] = 8'hD5;
mem[16'h2A0D] = 8'hAA;
mem[16'h2A0E] = 8'hD5;
mem[16'h2A0F] = 8'hAA;
mem[16'h2A10] = 8'hD5;
mem[16'h2A11] = 8'hAA;
mem[16'h2A12] = 8'hD5;
mem[16'h2A13] = 8'hAA;
mem[16'h2A14] = 8'hD5;
mem[16'h2A15] = 8'hAA;
mem[16'h2A16] = 8'hD5;
mem[16'h2A17] = 8'hAA;
mem[16'h2A18] = 8'hD5;
mem[16'h2A19] = 8'hAA;
mem[16'h2A1A] = 8'hD5;
mem[16'h2A1B] = 8'hAA;
mem[16'h2A1C] = 8'hD5;
mem[16'h2A1D] = 8'hAA;
mem[16'h2A1E] = 8'hD5;
mem[16'h2A1F] = 8'hAA;
mem[16'h2A20] = 8'hD5;
mem[16'h2A21] = 8'hAA;
mem[16'h2A22] = 8'hD5;
mem[16'h2A23] = 8'hAA;
mem[16'h2A24] = 8'h85;
mem[16'h2A25] = 8'h00;
mem[16'h2A26] = 8'h40;
mem[16'h2A27] = 8'h01;
mem[16'h2A28] = 8'h0A;
mem[16'h2A29] = 8'h51;
mem[16'h2A2A] = 8'h2A;
mem[16'h2A2B] = 8'h10;
mem[16'h2A2C] = 8'h28;
mem[16'h2A2D] = 8'h45;
mem[16'h2A2E] = 8'h2A;
mem[16'h2A2F] = 8'h51;
mem[16'h2A30] = 8'h0A;
mem[16'h2A31] = 8'h51;
mem[16'h2A32] = 8'h2A;
mem[16'h2A33] = 8'h10;
mem[16'h2A34] = 8'h28;
mem[16'h2A35] = 8'h45;
mem[16'h2A36] = 8'h2A;
mem[16'h2A37] = 8'h51;
mem[16'h2A38] = 8'h0A;
mem[16'h2A39] = 8'h51;
mem[16'h2A3A] = 8'h2A;
mem[16'h2A3B] = 8'h10;
mem[16'h2A3C] = 8'h28;
mem[16'h2A3D] = 8'h45;
mem[16'h2A3E] = 8'h2A;
mem[16'h2A3F] = 8'h51;
mem[16'h2A40] = 8'h0A;
mem[16'h2A41] = 8'h51;
mem[16'h2A42] = 8'h2A;
mem[16'h2A43] = 8'h10;
mem[16'h2A44] = 8'h28;
mem[16'h2A45] = 8'h45;
mem[16'h2A46] = 8'h2A;
mem[16'h2A47] = 8'h51;
mem[16'h2A48] = 8'h0A;
mem[16'h2A49] = 8'h51;
mem[16'h2A4A] = 8'h2A;
mem[16'h2A4B] = 8'h10;
mem[16'h2A4C] = 8'h08;
mem[16'h2A4D] = 8'h00;
mem[16'h2A4E] = 8'h00;
mem[16'h2A4F] = 8'h2A;
mem[16'h2A50] = 8'h00;
mem[16'h2A51] = 8'h00;
mem[16'h2A52] = 8'h00;
mem[16'h2A53] = 8'h00;
mem[16'h2A54] = 8'h00;
mem[16'h2A55] = 8'h00;
mem[16'h2A56] = 8'h00;
mem[16'h2A57] = 8'h00;
mem[16'h2A58] = 8'h00;
mem[16'h2A59] = 8'h00;
mem[16'h2A5A] = 8'h00;
mem[16'h2A5B] = 8'h00;
mem[16'h2A5C] = 8'h00;
mem[16'h2A5D] = 8'h00;
mem[16'h2A5E] = 8'h00;
mem[16'h2A5F] = 8'h00;
mem[16'h2A60] = 8'h00;
mem[16'h2A61] = 8'h00;
mem[16'h2A62] = 8'h00;
mem[16'h2A63] = 8'h00;
mem[16'h2A64] = 8'h00;
mem[16'h2A65] = 8'h00;
mem[16'h2A66] = 8'h00;
mem[16'h2A67] = 8'h00;
mem[16'h2A68] = 8'h00;
mem[16'h2A69] = 8'h00;
mem[16'h2A6A] = 8'h00;
mem[16'h2A6B] = 8'h00;
mem[16'h2A6C] = 8'h00;
mem[16'h2A6D] = 8'h00;
mem[16'h2A6E] = 8'h00;
mem[16'h2A6F] = 8'h00;
mem[16'h2A70] = 8'h00;
mem[16'h2A71] = 8'h00;
mem[16'h2A72] = 8'h00;
mem[16'h2A73] = 8'h00;
mem[16'h2A74] = 8'h00;
mem[16'h2A75] = 8'h00;
mem[16'h2A76] = 8'h00;
mem[16'h2A77] = 8'h2A;
mem[16'h2A78] = 8'h00;
mem[16'h2A79] = 8'h00;
mem[16'h2A7A] = 8'h00;
mem[16'h2A7B] = 8'h00;
mem[16'h2A7C] = 8'h00;
mem[16'h2A7D] = 8'h00;
mem[16'h2A7E] = 8'h00;
mem[16'h2A7F] = 8'h00;
mem[16'h2A80] = 8'hFD;
mem[16'h2A81] = 8'hD4;
mem[16'h2A82] = 8'hD2;
mem[16'h2A83] = 8'hCF;
mem[16'h2A84] = 8'hAA;
mem[16'h2A85] = 8'hAA;
mem[16'h2A86] = 8'hD5;
mem[16'h2A87] = 8'hAA;
mem[16'h2A88] = 8'hF5;
mem[16'h2A89] = 8'hD3;
mem[16'h2A8A] = 8'hCA;
mem[16'h2A8B] = 8'hBE;
mem[16'h2A8C] = 8'hAA;
mem[16'h2A8D] = 8'hA9;
mem[16'h2A8E] = 8'hD5;
mem[16'h2A8F] = 8'hAA;
mem[16'h2A90] = 8'hD5;
mem[16'h2A91] = 8'hCF;
mem[16'h2A92] = 8'hAA;
mem[16'h2A93] = 8'hFA;
mem[16'h2A94] = 8'hA9;
mem[16'h2A95] = 8'hA5;
mem[16'h2A96] = 8'hD5;
mem[16'h2A97] = 8'hAA;
mem[16'h2A98] = 8'hD5;
mem[16'h2A99] = 8'hBE;
mem[16'h2A9A] = 8'hAA;
mem[16'h2A9B] = 8'hE9;
mem[16'h2A9C] = 8'hA7;
mem[16'h2A9D] = 8'h95;
mem[16'h2A9E] = 8'hD5;
mem[16'h2A9F] = 8'hAA;
mem[16'h2AA0] = 8'hD5;
mem[16'h2AA1] = 8'hAA;
mem[16'h2AA2] = 8'hD5;
mem[16'h2AA3] = 8'hAA;
mem[16'h2AA4] = 8'h85;
mem[16'h2AA5] = 8'h00;
mem[16'h2AA6] = 8'h0E;
mem[16'h2AA7] = 8'h38;
mem[16'h2AA8] = 8'h00;
mem[16'h2AA9] = 8'h00;
mem[16'h2AAA] = 8'h00;
mem[16'h2AAB] = 8'h00;
mem[16'h2AAC] = 8'h00;
mem[16'h2AAD] = 8'h00;
mem[16'h2AAE] = 8'h00;
mem[16'h2AAF] = 8'h00;
mem[16'h2AB0] = 8'h00;
mem[16'h2AB1] = 8'h00;
mem[16'h2AB2] = 8'h00;
mem[16'h2AB3] = 8'h00;
mem[16'h2AB4] = 8'h00;
mem[16'h2AB5] = 8'h00;
mem[16'h2AB6] = 8'h00;
mem[16'h2AB7] = 8'h00;
mem[16'h2AB8] = 8'h00;
mem[16'h2AB9] = 8'h00;
mem[16'h2ABA] = 8'h00;
mem[16'h2ABB] = 8'h00;
mem[16'h2ABC] = 8'h00;
mem[16'h2ABD] = 8'h00;
mem[16'h2ABE] = 8'h00;
mem[16'h2ABF] = 8'h00;
mem[16'h2AC0] = 8'h00;
mem[16'h2AC1] = 8'h00;
mem[16'h2AC2] = 8'h00;
mem[16'h2AC3] = 8'h00;
mem[16'h2AC4] = 8'h00;
mem[16'h2AC5] = 8'h00;
mem[16'h2AC6] = 8'h00;
mem[16'h2AC7] = 8'h00;
mem[16'h2AC8] = 8'h00;
mem[16'h2AC9] = 8'h00;
mem[16'h2ACA] = 8'h00;
mem[16'h2ACB] = 8'h00;
mem[16'h2ACC] = 8'h00;
mem[16'h2ACD] = 8'h00;
mem[16'h2ACE] = 8'h00;
mem[16'h2ACF] = 8'h2A;
mem[16'h2AD0] = 8'h00;
mem[16'h2AD1] = 8'h00;
mem[16'h2AD2] = 8'h00;
mem[16'h2AD3] = 8'h00;
mem[16'h2AD4] = 8'h4F;
mem[16'h2AD5] = 8'h4A;
mem[16'h2AD6] = 8'h07;
mem[16'h2AD7] = 8'h00;
mem[16'h2AD8] = 8'h00;
mem[16'h2AD9] = 8'h00;
mem[16'h2ADA] = 8'h00;
mem[16'h2ADB] = 8'h00;
mem[16'h2ADC] = 8'h00;
mem[16'h2ADD] = 8'h00;
mem[16'h2ADE] = 8'h00;
mem[16'h2ADF] = 8'h00;
mem[16'h2AE0] = 8'h00;
mem[16'h2AE1] = 8'h00;
mem[16'h2AE2] = 8'h4F;
mem[16'h2AE3] = 8'h4A;
mem[16'h2AE4] = 8'h07;
mem[16'h2AE5] = 8'h00;
mem[16'h2AE6] = 8'h00;
mem[16'h2AE7] = 8'h00;
mem[16'h2AE8] = 8'h00;
mem[16'h2AE9] = 8'h00;
mem[16'h2AEA] = 8'h00;
mem[16'h2AEB] = 8'h00;
mem[16'h2AEC] = 8'h00;
mem[16'h2AED] = 8'h00;
mem[16'h2AEE] = 8'h00;
mem[16'h2AEF] = 8'h00;
mem[16'h2AF0] = 8'h4F;
mem[16'h2AF1] = 8'h4A;
mem[16'h2AF2] = 8'h07;
mem[16'h2AF3] = 8'h00;
mem[16'h2AF4] = 8'h00;
mem[16'h2AF5] = 8'h00;
mem[16'h2AF6] = 8'h00;
mem[16'h2AF7] = 8'h2A;
mem[16'h2AF8] = 8'h00;
mem[16'h2AF9] = 8'h00;
mem[16'h2AFA] = 8'h00;
mem[16'h2AFB] = 8'h00;
mem[16'h2AFC] = 8'h00;
mem[16'h2AFD] = 8'h00;
mem[16'h2AFE] = 8'h00;
mem[16'h2AFF] = 8'h00;
mem[16'h2B00] = 8'hD5;
mem[16'h2B01] = 8'hAA;
mem[16'h2B02] = 8'hD5;
mem[16'h2B03] = 8'hAA;
mem[16'h2B04] = 8'hD5;
mem[16'h2B05] = 8'hAA;
mem[16'h2B06] = 8'hD5;
mem[16'h2B07] = 8'hAA;
mem[16'h2B08] = 8'hD5;
mem[16'h2B09] = 8'hAA;
mem[16'h2B0A] = 8'hD5;
mem[16'h2B0B] = 8'hAA;
mem[16'h2B0C] = 8'hD5;
mem[16'h2B0D] = 8'hAA;
mem[16'h2B0E] = 8'hD5;
mem[16'h2B0F] = 8'hAA;
mem[16'h2B10] = 8'hD5;
mem[16'h2B11] = 8'hAA;
mem[16'h2B12] = 8'hD5;
mem[16'h2B13] = 8'hAA;
mem[16'h2B14] = 8'hD5;
mem[16'h2B15] = 8'hAA;
mem[16'h2B16] = 8'hD5;
mem[16'h2B17] = 8'hAA;
mem[16'h2B18] = 8'hD5;
mem[16'h2B19] = 8'hAA;
mem[16'h2B1A] = 8'hD5;
mem[16'h2B1B] = 8'hAA;
mem[16'h2B1C] = 8'hD5;
mem[16'h2B1D] = 8'hAA;
mem[16'h2B1E] = 8'hD5;
mem[16'h2B1F] = 8'hAA;
mem[16'h2B20] = 8'hD5;
mem[16'h2B21] = 8'hAA;
mem[16'h2B22] = 8'hD5;
mem[16'h2B23] = 8'hAA;
mem[16'h2B24] = 8'h85;
mem[16'h2B25] = 8'h00;
mem[16'h2B26] = 8'h70;
mem[16'h2B27] = 8'h07;
mem[16'h2B28] = 8'h00;
mem[16'h2B29] = 8'h00;
mem[16'h2B2A] = 8'h1E;
mem[16'h2B2B] = 8'h55;
mem[16'h2B2C] = 8'h0A;
mem[16'h2B2D] = 8'h00;
mem[16'h2B2E] = 8'h00;
mem[16'h2B2F] = 8'h00;
mem[16'h2B30] = 8'h00;
mem[16'h2B31] = 8'h00;
mem[16'h2B32] = 8'h00;
mem[16'h2B33] = 8'h00;
mem[16'h2B34] = 8'h00;
mem[16'h2B35] = 8'h00;
mem[16'h2B36] = 8'h00;
mem[16'h2B37] = 8'h00;
mem[16'h2B38] = 8'h1E;
mem[16'h2B39] = 8'h55;
mem[16'h2B3A] = 8'h0A;
mem[16'h2B3B] = 8'h00;
mem[16'h2B3C] = 8'h00;
mem[16'h2B3D] = 8'h00;
mem[16'h2B3E] = 8'h00;
mem[16'h2B3F] = 8'h00;
mem[16'h2B40] = 8'h00;
mem[16'h2B41] = 8'h00;
mem[16'h2B42] = 8'h00;
mem[16'h2B43] = 8'h00;
mem[16'h2B44] = 8'h00;
mem[16'h2B45] = 8'h00;
mem[16'h2B46] = 8'h00;
mem[16'h2B47] = 8'h00;
mem[16'h2B48] = 8'h00;
mem[16'h2B49] = 8'h00;
mem[16'h2B4A] = 8'h00;
mem[16'h2B4B] = 8'h00;
mem[16'h2B4C] = 8'h00;
mem[16'h2B4D] = 8'h00;
mem[16'h2B4E] = 8'h00;
mem[16'h2B4F] = 8'h2A;
mem[16'h2B50] = 8'h2A;
mem[16'h2B51] = 8'h45;
mem[16'h2B52] = 8'h2A;
mem[16'h2B53] = 8'h44;
mem[16'h2B54] = 8'h2A;
mem[16'h2B55] = 8'h41;
mem[16'h2B56] = 8'h20;
mem[16'h2B57] = 8'h15;
mem[16'h2B58] = 8'h2A;
mem[16'h2B59] = 8'h45;
mem[16'h2B5A] = 8'h2A;
mem[16'h2B5B] = 8'h44;
mem[16'h2B5C] = 8'h2A;
mem[16'h2B5D] = 8'h41;
mem[16'h2B5E] = 8'h20;
mem[16'h2B5F] = 8'h15;
mem[16'h2B60] = 8'h2A;
mem[16'h2B61] = 8'h45;
mem[16'h2B62] = 8'h60;
mem[16'h2B63] = 8'h03;
mem[16'h2B64] = 8'h2A;
mem[16'h2B65] = 8'h41;
mem[16'h2B66] = 8'h20;
mem[16'h2B67] = 8'h15;
mem[16'h2B68] = 8'h2A;
mem[16'h2B69] = 8'h45;
mem[16'h2B6A] = 8'h2A;
mem[16'h2B6B] = 8'h44;
mem[16'h2B6C] = 8'h2A;
mem[16'h2B6D] = 8'h41;
mem[16'h2B6E] = 8'h20;
mem[16'h2B6F] = 8'h15;
mem[16'h2B70] = 8'h2A;
mem[16'h2B71] = 8'h45;
mem[16'h2B72] = 8'h2A;
mem[16'h2B73] = 8'h44;
mem[16'h2B74] = 8'h0A;
mem[16'h2B75] = 8'h00;
mem[16'h2B76] = 8'h00;
mem[16'h2B77] = 8'h2A;
mem[16'h2B78] = 8'h00;
mem[16'h2B79] = 8'h00;
mem[16'h2B7A] = 8'h00;
mem[16'h2B7B] = 8'h00;
mem[16'h2B7C] = 8'h00;
mem[16'h2B7D] = 8'h00;
mem[16'h2B7E] = 8'h00;
mem[16'h2B7F] = 8'h00;
mem[16'h2B80] = 8'hAB;
mem[16'h2B81] = 8'hAB;
mem[16'h2B82] = 8'hD5;
mem[16'h2B83] = 8'hAA;
mem[16'h2B84] = 8'hD5;
mem[16'h2B85] = 8'hAA;
mem[16'h2B86] = 8'hD5;
mem[16'h2B87] = 8'hAA;
mem[16'h2B88] = 8'hD5;
mem[16'h2B89] = 8'hAA;
mem[16'h2B8A] = 8'hD5;
mem[16'h2B8B] = 8'hD6;
mem[16'h2B8C] = 8'hAA;
mem[16'h2B8D] = 8'hD5;
mem[16'h2B8E] = 8'hAA;
mem[16'h2B8F] = 8'hD5;
mem[16'h2B90] = 8'hAA;
mem[16'h2B91] = 8'hD5;
mem[16'h2B92] = 8'hAA;
mem[16'h2B93] = 8'hD5;
mem[16'h2B94] = 8'hAA;
mem[16'h2B95] = 8'hD5;
mem[16'h2B96] = 8'hAA;
mem[16'h2B97] = 8'hD5;
mem[16'h2B98] = 8'hAA;
mem[16'h2B99] = 8'hB5;
mem[16'h2B9A] = 8'hD5;
mem[16'h2B9B] = 8'hAA;
mem[16'h2B9C] = 8'hD5;
mem[16'h2B9D] = 8'hAA;
mem[16'h2B9E] = 8'hD5;
mem[16'h2B9F] = 8'hAA;
mem[16'h2BA0] = 8'hD5;
mem[16'h2BA1] = 8'hAA;
mem[16'h2BA2] = 8'hD5;
mem[16'h2BA3] = 8'hAA;
mem[16'h2BA4] = 8'h85;
mem[16'h2BA5] = 8'h00;
mem[16'h2BA6] = 8'h00;
mem[16'h2BA7] = 8'h00;
mem[16'h2BA8] = 8'h00;
mem[16'h2BA9] = 8'hF0;
mem[16'h2BAA] = 8'hC0;
mem[16'h2BAB] = 8'h83;
mem[16'h2BAC] = 8'h00;
mem[16'h2BAD] = 8'h00;
mem[16'h2BAE] = 8'h00;
mem[16'h2BAF] = 8'h00;
mem[16'h2BB0] = 8'h00;
mem[16'h2BB1] = 8'h00;
mem[16'h2BB2] = 8'h00;
mem[16'h2BB3] = 8'h00;
mem[16'h2BB4] = 8'h00;
mem[16'h2BB5] = 8'h00;
mem[16'h2BB6] = 8'h00;
mem[16'h2BB7] = 8'h00;
mem[16'h2BB8] = 8'h00;
mem[16'h2BB9] = 8'h00;
mem[16'h2BBA] = 8'h00;
mem[16'h2BBB] = 8'h00;
mem[16'h2BBC] = 8'h00;
mem[16'h2BBD] = 8'h00;
mem[16'h2BBE] = 8'h00;
mem[16'h2BBF] = 8'h00;
mem[16'h2BC0] = 8'h00;
mem[16'h2BC1] = 8'h00;
mem[16'h2BC2] = 8'h00;
mem[16'h2BC3] = 8'h00;
mem[16'h2BC4] = 8'h00;
mem[16'h2BC5] = 8'h00;
mem[16'h2BC6] = 8'h00;
mem[16'h2BC7] = 8'h00;
mem[16'h2BC8] = 8'h00;
mem[16'h2BC9] = 8'h00;
mem[16'h2BCA] = 8'h00;
mem[16'h2BCB] = 8'h00;
mem[16'h2BCC] = 8'h00;
mem[16'h2BCD] = 8'h00;
mem[16'h2BCE] = 8'h00;
mem[16'h2BCF] = 8'h2A;
mem[16'h2BD0] = 8'h2A;
mem[16'h2BD1] = 8'h45;
mem[16'h2BD2] = 8'h2A;
mem[16'h2BD3] = 8'h44;
mem[16'h2BD4] = 8'h2A;
mem[16'h2BD5] = 8'h41;
mem[16'h2BD6] = 8'h20;
mem[16'h2BD7] = 8'h15;
mem[16'h2BD8] = 8'h2A;
mem[16'h2BD9] = 8'h45;
mem[16'h2BDA] = 8'h2A;
mem[16'h2BDB] = 8'h44;
mem[16'h2BDC] = 8'h2A;
mem[16'h2BDD] = 8'h41;
mem[16'h2BDE] = 8'h20;
mem[16'h2BDF] = 8'h15;
mem[16'h2BE0] = 8'h2A;
mem[16'h2BE1] = 8'h45;
mem[16'h2BE2] = 8'h0E;
mem[16'h2BE3] = 8'h38;
mem[16'h2BE4] = 8'h2A;
mem[16'h2BE5] = 8'h41;
mem[16'h2BE6] = 8'h20;
mem[16'h2BE7] = 8'h15;
mem[16'h2BE8] = 8'h2A;
mem[16'h2BE9] = 8'h45;
mem[16'h2BEA] = 8'h2A;
mem[16'h2BEB] = 8'h44;
mem[16'h2BEC] = 8'h2A;
mem[16'h2BED] = 8'h41;
mem[16'h2BEE] = 8'h20;
mem[16'h2BEF] = 8'h15;
mem[16'h2BF0] = 8'h2A;
mem[16'h2BF1] = 8'h45;
mem[16'h2BF2] = 8'h2A;
mem[16'h2BF3] = 8'h44;
mem[16'h2BF4] = 8'h0A;
mem[16'h2BF5] = 8'h4A;
mem[16'h2BF6] = 8'h00;
mem[16'h2BF7] = 8'h2A;
mem[16'h2BF8] = 8'h00;
mem[16'h2BF9] = 8'h00;
mem[16'h2BFA] = 8'h00;
mem[16'h2BFB] = 8'h00;
mem[16'h2BFC] = 8'h00;
mem[16'h2BFD] = 8'h00;
mem[16'h2BFE] = 8'h00;
mem[16'h2BFF] = 8'h00;
mem[16'h2C00] = 8'h00;
mem[16'h2C01] = 8'h7E;
mem[16'h2C02] = 8'h10;
mem[16'h2C03] = 8'h00;
mem[16'h2C04] = 8'h3C;
mem[16'h2C05] = 8'h02;
mem[16'h2C06] = 8'h44;
mem[16'h2C07] = 8'h46;
mem[16'h2C08] = 8'h42;
mem[16'h2C09] = 8'h00;
mem[16'h2C0A] = 8'h42;
mem[16'h2C0B] = 8'h42;
mem[16'h2C0C] = 8'h42;
mem[16'h2C0D] = 8'h42;
mem[16'h2C0E] = 8'h42;
mem[16'h2C0F] = 8'h42;
mem[16'h2C10] = 8'h00;
mem[16'h2C11] = 8'h00;
mem[16'h2C12] = 8'h00;
mem[16'h2C13] = 8'h00;
mem[16'h2C14] = 8'h38;
mem[16'h2C15] = 8'h44;
mem[16'h2C16] = 8'h42;
mem[16'h2C17] = 8'h46;
mem[16'h2C18] = 8'h00;
mem[16'h2C19] = 8'h3C;
mem[16'h2C1A] = 8'h02;
mem[16'h2C1B] = 8'h44;
mem[16'h2C1C] = 8'h46;
mem[16'h2C1D] = 8'h42;
mem[16'h2C1E] = 8'h00;
mem[16'h2C1F] = 8'h42;
mem[16'h2C20] = 8'h42;
mem[16'h2C21] = 8'h42;
mem[16'h2C22] = 8'h42;
mem[16'h2C23] = 8'h42;
mem[16'h2C24] = 8'h42;
mem[16'h2C25] = 8'h00;
mem[16'h2C26] = 8'h40;
mem[16'h2C27] = 8'h01;
mem[16'h2C28] = 8'hD5;
mem[16'h2C29] = 8'hAA;
mem[16'h2C2A] = 8'hD5;
mem[16'h2C2B] = 8'hAA;
mem[16'h2C2C] = 8'hB5;
mem[16'h2C2D] = 8'hD5;
mem[16'h2C2E] = 8'hAA;
mem[16'h2C2F] = 8'hD5;
mem[16'h2C30] = 8'hAA;
mem[16'h2C31] = 8'hD5;
mem[16'h2C32] = 8'hAA;
mem[16'h2C33] = 8'hD5;
mem[16'h2C34] = 8'hD6;
mem[16'h2C35] = 8'hAA;
mem[16'h2C36] = 8'hD5;
mem[16'h2C37] = 8'hAA;
mem[16'h2C38] = 8'hD5;
mem[16'h2C39] = 8'hD5;
mem[16'h2C3A] = 8'hAA;
mem[16'h2C3B] = 8'hD5;
mem[16'h2C3C] = 8'hAA;
mem[16'h2C3D] = 8'hD5;
mem[16'h2C3E] = 8'hAA;
mem[16'h2C3F] = 8'hD5;
mem[16'h2C40] = 8'hDA;
mem[16'h2C41] = 8'hAA;
mem[16'h2C42] = 8'hD5;
mem[16'h2C43] = 8'hAA;
mem[16'h2C44] = 8'hAB;
mem[16'h2C45] = 8'hD5;
mem[16'h2C46] = 8'hAA;
mem[16'h2C47] = 8'hD5;
mem[16'h2C48] = 8'hAA;
mem[16'h2C49] = 8'hD5;
mem[16'h2C4A] = 8'hAA;
mem[16'h2C4B] = 8'hB5;
mem[16'h2C4C] = 8'h85;
mem[16'h2C4D] = 8'h00;
mem[16'h2C4E] = 8'h00;
mem[16'h2C4F] = 8'h00;
mem[16'h2C50] = 8'h00;
mem[16'h2C51] = 8'h00;
mem[16'h2C52] = 8'h00;
mem[16'h2C53] = 8'h00;
mem[16'h2C54] = 8'h00;
mem[16'h2C55] = 8'h00;
mem[16'h2C56] = 8'h00;
mem[16'h2C57] = 8'h00;
mem[16'h2C58] = 8'h00;
mem[16'h2C59] = 8'h00;
mem[16'h2C5A] = 8'h00;
mem[16'h2C5B] = 8'h00;
mem[16'h2C5C] = 8'h00;
mem[16'h2C5D] = 8'h00;
mem[16'h2C5E] = 8'h00;
mem[16'h2C5F] = 8'h00;
mem[16'h2C60] = 8'h00;
mem[16'h2C61] = 8'h00;
mem[16'h2C62] = 8'h00;
mem[16'h2C63] = 8'h00;
mem[16'h2C64] = 8'h00;
mem[16'h2C65] = 8'h00;
mem[16'h2C66] = 8'h00;
mem[16'h2C67] = 8'h00;
mem[16'h2C68] = 8'h00;
mem[16'h2C69] = 8'h00;
mem[16'h2C6A] = 8'h00;
mem[16'h2C6B] = 8'h00;
mem[16'h2C6C] = 8'h00;
mem[16'h2C6D] = 8'h00;
mem[16'h2C6E] = 8'h00;
mem[16'h2C6F] = 8'h00;
mem[16'h2C70] = 8'h00;
mem[16'h2C71] = 8'h00;
mem[16'h2C72] = 8'h00;
mem[16'h2C73] = 8'h00;
mem[16'h2C74] = 8'h00;
mem[16'h2C75] = 8'h00;
mem[16'h2C76] = 8'h00;
mem[16'h2C77] = 8'h2A;
mem[16'h2C78] = 8'h00;
mem[16'h2C79] = 8'h00;
mem[16'h2C7A] = 8'h00;
mem[16'h2C7B] = 8'h00;
mem[16'h2C7C] = 8'h00;
mem[16'h2C7D] = 8'h00;
mem[16'h2C7E] = 8'h00;
mem[16'h2C7F] = 8'h00;
mem[16'h2C80] = 8'h28;
mem[16'h2C81] = 8'h15;
mem[16'h2C82] = 8'h08;
mem[16'h2C83] = 8'hAA;
mem[16'h2C84] = 8'hD5;
mem[16'h2C85] = 8'h55;
mem[16'h2C86] = 8'h28;
mem[16'h2C87] = 8'h45;
mem[16'h2C88] = 8'h28;
mem[16'h2C89] = 8'h15;
mem[16'h2C8A] = 8'hD5;
mem[16'h2C8B] = 8'hAA;
mem[16'h2C8C] = 8'h22;
mem[16'h2C8D] = 8'h55;
mem[16'h2C8E] = 8'h28;
mem[16'h2C8F] = 8'h45;
mem[16'h2C90] = 8'hD5;
mem[16'h2C91] = 8'hAA;
mem[16'h2C92] = 8'h08;
mem[16'h2C93] = 8'h54;
mem[16'h2C94] = 8'h22;
mem[16'h2C95] = 8'h55;
mem[16'h2C96] = 8'h28;
mem[16'h2C97] = 8'hAA;
mem[16'h2C98] = 8'hD5;
mem[16'h2C99] = 8'h15;
mem[16'h2C9A] = 8'h08;
mem[16'h2C9B] = 8'h54;
mem[16'h2C9C] = 8'h22;
mem[16'h2C9D] = 8'hAA;
mem[16'h2C9E] = 8'hD5;
mem[16'h2C9F] = 8'h45;
mem[16'h2CA0] = 8'h28;
mem[16'h2CA1] = 8'h15;
mem[16'h2CA2] = 8'h08;
mem[16'h2CA3] = 8'h54;
mem[16'h2CA4] = 8'h02;
mem[16'h2CA5] = 8'h00;
mem[16'h2CA6] = 8'h7C;
mem[16'h2CA7] = 8'h1F;
mem[16'h2CA8] = 8'hD5;
mem[16'h2CA9] = 8'hAA;
mem[16'h2CAA] = 8'hD5;
mem[16'h2CAB] = 8'hAA;
mem[16'h2CAC] = 8'hD5;
mem[16'h2CAD] = 8'hAA;
mem[16'h2CAE] = 8'hD5;
mem[16'h2CAF] = 8'hAA;
mem[16'h2CB0] = 8'hD5;
mem[16'h2CB1] = 8'hAA;
mem[16'h2CB2] = 8'hD5;
mem[16'h2CB3] = 8'hAA;
mem[16'h2CB4] = 8'hD5;
mem[16'h2CB5] = 8'hAA;
mem[16'h2CB6] = 8'hD5;
mem[16'h2CB7] = 8'hAA;
mem[16'h2CB8] = 8'hD5;
mem[16'h2CB9] = 8'hAA;
mem[16'h2CBA] = 8'hD5;
mem[16'h2CBB] = 8'hAA;
mem[16'h2CBC] = 8'hD5;
mem[16'h2CBD] = 8'hAA;
mem[16'h2CBE] = 8'hD5;
mem[16'h2CBF] = 8'hAA;
mem[16'h2CC0] = 8'hD5;
mem[16'h2CC1] = 8'hAA;
mem[16'h2CC2] = 8'hD5;
mem[16'h2CC3] = 8'hAA;
mem[16'h2CC4] = 8'hD5;
mem[16'h2CC5] = 8'hAA;
mem[16'h2CC6] = 8'hD5;
mem[16'h2CC7] = 8'hAA;
mem[16'h2CC8] = 8'hD5;
mem[16'h2CC9] = 8'hAA;
mem[16'h2CCA] = 8'hD5;
mem[16'h2CCB] = 8'hAA;
mem[16'h2CCC] = 8'h85;
mem[16'h2CCD] = 8'h00;
mem[16'h2CCE] = 8'h00;
mem[16'h2CCF] = 8'h2A;
mem[16'h2CD0] = 8'h00;
mem[16'h2CD1] = 8'h00;
mem[16'h2CD2] = 8'h00;
mem[16'h2CD3] = 8'h00;
mem[16'h2CD4] = 8'h00;
mem[16'h2CD5] = 8'h55;
mem[16'h2CD6] = 8'h28;
mem[16'h2CD7] = 8'h03;
mem[16'h2CD8] = 8'h00;
mem[16'h2CD9] = 8'h00;
mem[16'h2CDA] = 8'h00;
mem[16'h2CDB] = 8'h00;
mem[16'h2CDC] = 8'h00;
mem[16'h2CDD] = 8'h00;
mem[16'h2CDE] = 8'h00;
mem[16'h2CDF] = 8'h00;
mem[16'h2CE0] = 8'h00;
mem[16'h2CE1] = 8'h55;
mem[16'h2CE2] = 8'h28;
mem[16'h2CE3] = 8'h03;
mem[16'h2CE4] = 8'h00;
mem[16'h2CE5] = 8'h00;
mem[16'h2CE6] = 8'h00;
mem[16'h2CE7] = 8'h00;
mem[16'h2CE8] = 8'h00;
mem[16'h2CE9] = 8'h00;
mem[16'h2CEA] = 8'h00;
mem[16'h2CEB] = 8'h00;
mem[16'h2CEC] = 8'h00;
mem[16'h2CED] = 8'h55;
mem[16'h2CEE] = 8'h28;
mem[16'h2CEF] = 8'h03;
mem[16'h2CF0] = 8'h00;
mem[16'h2CF1] = 8'h00;
mem[16'h2CF2] = 8'h00;
mem[16'h2CF3] = 8'h00;
mem[16'h2CF4] = 8'h00;
mem[16'h2CF5] = 8'h00;
mem[16'h2CF6] = 8'h00;
mem[16'h2CF7] = 8'h2A;
mem[16'h2CF8] = 8'h00;
mem[16'h2CF9] = 8'h00;
mem[16'h2CFA] = 8'h00;
mem[16'h2CFB] = 8'h00;
mem[16'h2CFC] = 8'h00;
mem[16'h2CFD] = 8'h00;
mem[16'h2CFE] = 8'h00;
mem[16'h2CFF] = 8'h00;
mem[16'h2D00] = 8'h28;
mem[16'h2D01] = 8'h15;
mem[16'h2D02] = 8'h08;
mem[16'h2D03] = 8'hAA;
mem[16'h2D04] = 8'hD5;
mem[16'h2D05] = 8'h55;
mem[16'h2D06] = 8'h28;
mem[16'h2D07] = 8'h45;
mem[16'h2D08] = 8'h28;
mem[16'h2D09] = 8'h15;
mem[16'h2D0A] = 8'hD5;
mem[16'h2D0B] = 8'hAA;
mem[16'h2D0C] = 8'h22;
mem[16'h2D0D] = 8'h55;
mem[16'h2D0E] = 8'h28;
mem[16'h2D0F] = 8'h45;
mem[16'h2D10] = 8'hD5;
mem[16'h2D11] = 8'hAA;
mem[16'h2D12] = 8'h08;
mem[16'h2D13] = 8'h54;
mem[16'h2D14] = 8'h22;
mem[16'h2D15] = 8'h55;
mem[16'h2D16] = 8'h28;
mem[16'h2D17] = 8'hAA;
mem[16'h2D18] = 8'hD5;
mem[16'h2D19] = 8'h15;
mem[16'h2D1A] = 8'h08;
mem[16'h2D1B] = 8'h54;
mem[16'h2D1C] = 8'h22;
mem[16'h2D1D] = 8'hAA;
mem[16'h2D1E] = 8'hD5;
mem[16'h2D1F] = 8'h45;
mem[16'h2D20] = 8'h28;
mem[16'h2D21] = 8'h15;
mem[16'h2D22] = 8'h08;
mem[16'h2D23] = 8'h54;
mem[16'h2D24] = 8'h02;
mem[16'h2D25] = 8'h00;
mem[16'h2D26] = 8'h60;
mem[16'h2D27] = 8'h03;
mem[16'h2D28] = 8'hD5;
mem[16'h2D29] = 8'hAA;
mem[16'h2D2A] = 8'hD5;
mem[16'h2D2B] = 8'hAA;
mem[16'h2D2C] = 8'hD5;
mem[16'h2D2D] = 8'hD6;
mem[16'h2D2E] = 8'hCA;
mem[16'h2D2F] = 8'hEA;
mem[16'h2D30] = 8'hAA;
mem[16'h2D31] = 8'hA9;
mem[16'h2D32] = 8'hAD;
mem[16'h2D33] = 8'h95;
mem[16'h2D34] = 8'hD5;
mem[16'h2D35] = 8'hAA;
mem[16'h2D36] = 8'hD5;
mem[16'h2D37] = 8'hAA;
mem[16'h2D38] = 8'hD5;
mem[16'h2D39] = 8'hAA;
mem[16'h2D3A] = 8'hD5;
mem[16'h2D3B] = 8'hAA;
mem[16'h2D3C] = 8'hAB;
mem[16'h2D3D] = 8'hA5;
mem[16'h2D3E] = 8'hB5;
mem[16'h2D3F] = 8'hD5;
mem[16'h2D40] = 8'hD4;
mem[16'h2D41] = 8'hD6;
mem[16'h2D42] = 8'hCA;
mem[16'h2D43] = 8'hAA;
mem[16'h2D44] = 8'hD5;
mem[16'h2D45] = 8'hAA;
mem[16'h2D46] = 8'hD5;
mem[16'h2D47] = 8'hAA;
mem[16'h2D48] = 8'hD5;
mem[16'h2D49] = 8'hAA;
mem[16'h2D4A] = 8'hD5;
mem[16'h2D4B] = 8'hAA;
mem[16'h2D4C] = 8'h85;
mem[16'h2D4D] = 8'h00;
mem[16'h2D4E] = 8'h00;
mem[16'h2D4F] = 8'h2A;
mem[16'h2D50] = 8'h00;
mem[16'h2D51] = 8'h00;
mem[16'h2D52] = 8'h00;
mem[16'h2D53] = 8'h00;
mem[16'h2D54] = 8'h00;
mem[16'h2D55] = 8'h00;
mem[16'h2D56] = 8'h00;
mem[16'h2D57] = 8'h00;
mem[16'h2D58] = 8'h00;
mem[16'h2D59] = 8'h00;
mem[16'h2D5A] = 8'h00;
mem[16'h2D5B] = 8'h00;
mem[16'h2D5C] = 8'h00;
mem[16'h2D5D] = 8'h00;
mem[16'h2D5E] = 8'h00;
mem[16'h2D5F] = 8'h00;
mem[16'h2D60] = 8'h00;
mem[16'h2D61] = 8'h00;
mem[16'h2D62] = 8'h00;
mem[16'h2D63] = 8'h00;
mem[16'h2D64] = 8'h00;
mem[16'h2D65] = 8'h00;
mem[16'h2D66] = 8'h00;
mem[16'h2D67] = 8'h00;
mem[16'h2D68] = 8'h00;
mem[16'h2D69] = 8'h00;
mem[16'h2D6A] = 8'h00;
mem[16'h2D6B] = 8'h00;
mem[16'h2D6C] = 8'h00;
mem[16'h2D6D] = 8'h00;
mem[16'h2D6E] = 8'h00;
mem[16'h2D6F] = 8'h00;
mem[16'h2D70] = 8'h00;
mem[16'h2D71] = 8'h00;
mem[16'h2D72] = 8'h00;
mem[16'h2D73] = 8'h00;
mem[16'h2D74] = 8'h00;
mem[16'h2D75] = 8'h00;
mem[16'h2D76] = 8'h00;
mem[16'h2D77] = 8'h2A;
mem[16'h2D78] = 8'h00;
mem[16'h2D79] = 8'h00;
mem[16'h2D7A] = 8'h00;
mem[16'h2D7B] = 8'h00;
mem[16'h2D7C] = 8'h00;
mem[16'h2D7D] = 8'h00;
mem[16'h2D7E] = 8'h00;
mem[16'h2D7F] = 8'h00;
mem[16'h2D80] = 8'hD5;
mem[16'h2D81] = 8'hAA;
mem[16'h2D82] = 8'hD5;
mem[16'h2D83] = 8'hAA;
mem[16'h2D84] = 8'hD5;
mem[16'h2D85] = 8'hAA;
mem[16'h2D86] = 8'hAB;
mem[16'h2D87] = 8'hD5;
mem[16'h2D88] = 8'hAA;
mem[16'h2D89] = 8'hD5;
mem[16'h2D8A] = 8'hAA;
mem[16'h2D8B] = 8'hD5;
mem[16'h2D8C] = 8'hAA;
mem[16'h2D8D] = 8'hD5;
mem[16'h2D8E] = 8'hAA;
mem[16'h2D8F] = 8'hD5;
mem[16'h2D90] = 8'hD5;
mem[16'h2D91] = 8'hAA;
mem[16'h2D92] = 8'hAD;
mem[16'h2D93] = 8'hD5;
mem[16'h2D94] = 8'hAA;
mem[16'h2D95] = 8'hD5;
mem[16'h2D96] = 8'hAA;
mem[16'h2D97] = 8'hD5;
mem[16'h2D98] = 8'hAA;
mem[16'h2D99] = 8'hD5;
mem[16'h2D9A] = 8'hAA;
mem[16'h2D9B] = 8'hD5;
mem[16'h2D9C] = 8'hD6;
mem[16'h2D9D] = 8'hAA;
mem[16'h2D9E] = 8'hD5;
mem[16'h2D9F] = 8'hAA;
mem[16'h2DA0] = 8'hD5;
mem[16'h2DA1] = 8'hAA;
mem[16'h2DA2] = 8'hD5;
mem[16'h2DA3] = 8'hAA;
mem[16'h2DA4] = 8'h85;
mem[16'h2DA5] = 8'h00;
mem[16'h2DA6] = 8'h0E;
mem[16'h2DA7] = 8'h38;
mem[16'h2DA8] = 8'h0A;
mem[16'h2DA9] = 8'h04;
mem[16'h2DAA] = 8'h2A;
mem[16'h2DAB] = 8'h51;
mem[16'h2DAC] = 8'h2A;
mem[16'h2DAD] = 8'h54;
mem[16'h2DAE] = 8'h22;
mem[16'h2DAF] = 8'h54;
mem[16'h2DB0] = 8'h0A;
mem[16'h2DB1] = 8'h04;
mem[16'h2DB2] = 8'h2A;
mem[16'h2DB3] = 8'h51;
mem[16'h2DB4] = 8'h2A;
mem[16'h2DB5] = 8'h54;
mem[16'h2DB6] = 8'h22;
mem[16'h2DB7] = 8'h54;
mem[16'h2DB8] = 8'h0A;
mem[16'h2DB9] = 8'h04;
mem[16'h2DBA] = 8'h2A;
mem[16'h2DBB] = 8'h51;
mem[16'h2DBC] = 8'h2A;
mem[16'h2DBD] = 8'h54;
mem[16'h2DBE] = 8'h22;
mem[16'h2DBF] = 8'h54;
mem[16'h2DC0] = 8'h0A;
mem[16'h2DC1] = 8'h04;
mem[16'h2DC2] = 8'h2A;
mem[16'h2DC3] = 8'h51;
mem[16'h2DC4] = 8'h2A;
mem[16'h2DC5] = 8'h54;
mem[16'h2DC6] = 8'h22;
mem[16'h2DC7] = 8'h54;
mem[16'h2DC8] = 8'h0A;
mem[16'h2DC9] = 8'h04;
mem[16'h2DCA] = 8'h2A;
mem[16'h2DCB] = 8'h51;
mem[16'h2DCC] = 8'h0A;
mem[16'h2DCD] = 8'h00;
mem[16'h2DCE] = 8'h00;
mem[16'h2DCF] = 8'h2A;
mem[16'h2DD0] = 8'h00;
mem[16'h2DD1] = 8'hA8;
mem[16'h2DD2] = 8'h95;
mem[16'h2DD3] = 8'h81;
mem[16'h2DD4] = 8'h00;
mem[16'h2DD5] = 8'h00;
mem[16'h2DD6] = 8'h00;
mem[16'h2DD7] = 8'h00;
mem[16'h2DD8] = 8'h00;
mem[16'h2DD9] = 8'h00;
mem[16'h2DDA] = 8'h00;
mem[16'h2DDB] = 8'hC0;
mem[16'h2DDC] = 8'hAA;
mem[16'h2DDD] = 8'h89;
mem[16'h2DDE] = 8'h00;
mem[16'h2DDF] = 8'h00;
mem[16'h2DE0] = 8'h00;
mem[16'h2DE1] = 8'h00;
mem[16'h2DE2] = 8'h00;
mem[16'h2DE3] = 8'h00;
mem[16'h2DE4] = 8'h00;
mem[16'h2DE5] = 8'h00;
mem[16'h2DE6] = 8'hD4;
mem[16'h2DE7] = 8'hCA;
mem[16'h2DE8] = 8'h80;
mem[16'h2DE9] = 8'h00;
mem[16'h2DEA] = 8'h00;
mem[16'h2DEB] = 8'h00;
mem[16'h2DEC] = 8'h00;
mem[16'h2DED] = 8'h00;
mem[16'h2DEE] = 8'h00;
mem[16'h2DEF] = 8'h00;
mem[16'h2DF0] = 8'h00;
mem[16'h2DF1] = 8'h00;
mem[16'h2DF2] = 8'h00;
mem[16'h2DF3] = 8'h00;
mem[16'h2DF4] = 8'h00;
mem[16'h2DF5] = 8'h00;
mem[16'h2DF6] = 8'h00;
mem[16'h2DF7] = 8'h2A;
mem[16'h2DF8] = 8'h00;
mem[16'h2DF9] = 8'h00;
mem[16'h2DFA] = 8'h00;
mem[16'h2DFB] = 8'h00;
mem[16'h2DFC] = 8'h00;
mem[16'h2DFD] = 8'h00;
mem[16'h2DFE] = 8'h00;
mem[16'h2DFF] = 8'h00;
mem[16'h2E00] = 8'hD5;
mem[16'h2E01] = 8'hAA;
mem[16'h2E02] = 8'hD5;
mem[16'h2E03] = 8'hAA;
mem[16'h2E04] = 8'hD5;
mem[16'h2E05] = 8'hAA;
mem[16'h2E06] = 8'hD5;
mem[16'h2E07] = 8'hAA;
mem[16'h2E08] = 8'hD5;
mem[16'h2E09] = 8'hAA;
mem[16'h2E0A] = 8'hD5;
mem[16'h2E0B] = 8'hAA;
mem[16'h2E0C] = 8'hD5;
mem[16'h2E0D] = 8'hAA;
mem[16'h2E0E] = 8'hD5;
mem[16'h2E0F] = 8'hAA;
mem[16'h2E10] = 8'hD5;
mem[16'h2E11] = 8'hAA;
mem[16'h2E12] = 8'hD5;
mem[16'h2E13] = 8'hAA;
mem[16'h2E14] = 8'hD5;
mem[16'h2E15] = 8'hAA;
mem[16'h2E16] = 8'hD5;
mem[16'h2E17] = 8'hAA;
mem[16'h2E18] = 8'hD5;
mem[16'h2E19] = 8'hAA;
mem[16'h2E1A] = 8'hD5;
mem[16'h2E1B] = 8'hAA;
mem[16'h2E1C] = 8'hD5;
mem[16'h2E1D] = 8'hAA;
mem[16'h2E1E] = 8'hD5;
mem[16'h2E1F] = 8'hAA;
mem[16'h2E20] = 8'hD5;
mem[16'h2E21] = 8'hAA;
mem[16'h2E22] = 8'hD5;
mem[16'h2E23] = 8'hAA;
mem[16'h2E24] = 8'h85;
mem[16'h2E25] = 8'h00;
mem[16'h2E26] = 8'h60;
mem[16'h2E27] = 8'h03;
mem[16'h2E28] = 8'h2A;
mem[16'h2E29] = 8'h54;
mem[16'h2E2A] = 8'h0A;
mem[16'h2E2B] = 8'h55;
mem[16'h2E2C] = 8'h08;
mem[16'h2E2D] = 8'h55;
mem[16'h2E2E] = 8'h02;
mem[16'h2E2F] = 8'h41;
mem[16'h2E30] = 8'h2A;
mem[16'h2E31] = 8'h54;
mem[16'h2E32] = 8'h0A;
mem[16'h2E33] = 8'h55;
mem[16'h2E34] = 8'h08;
mem[16'h2E35] = 8'h55;
mem[16'h2E36] = 8'h02;
mem[16'h2E37] = 8'h41;
mem[16'h2E38] = 8'h2A;
mem[16'h2E39] = 8'h54;
mem[16'h2E3A] = 8'h0A;
mem[16'h2E3B] = 8'h55;
mem[16'h2E3C] = 8'h08;
mem[16'h2E3D] = 8'h55;
mem[16'h2E3E] = 8'h02;
mem[16'h2E3F] = 8'h41;
mem[16'h2E40] = 8'h2A;
mem[16'h2E41] = 8'h54;
mem[16'h2E42] = 8'h0A;
mem[16'h2E43] = 8'h55;
mem[16'h2E44] = 8'h08;
mem[16'h2E45] = 8'h55;
mem[16'h2E46] = 8'h02;
mem[16'h2E47] = 8'h41;
mem[16'h2E48] = 8'h2A;
mem[16'h2E49] = 8'h54;
mem[16'h2E4A] = 8'h0A;
mem[16'h2E4B] = 8'h55;
mem[16'h2E4C] = 8'h08;
mem[16'h2E4D] = 8'h00;
mem[16'h2E4E] = 8'h00;
mem[16'h2E4F] = 8'h2A;
mem[16'h2E50] = 8'h00;
mem[16'h2E51] = 8'h00;
mem[16'h2E52] = 8'h00;
mem[16'h2E53] = 8'h00;
mem[16'h2E54] = 8'h0F;
mem[16'h2E55] = 8'h40;
mem[16'h2E56] = 8'h07;
mem[16'h2E57] = 8'h00;
mem[16'h2E58] = 8'h00;
mem[16'h2E59] = 8'h00;
mem[16'h2E5A] = 8'h00;
mem[16'h2E5B] = 8'h00;
mem[16'h2E5C] = 8'h00;
mem[16'h2E5D] = 8'h00;
mem[16'h2E5E] = 8'h00;
mem[16'h2E5F] = 8'h00;
mem[16'h2E60] = 8'h00;
mem[16'h2E61] = 8'h00;
mem[16'h2E62] = 8'h0F;
mem[16'h2E63] = 8'h40;
mem[16'h2E64] = 8'h07;
mem[16'h2E65] = 8'h00;
mem[16'h2E66] = 8'h00;
mem[16'h2E67] = 8'h00;
mem[16'h2E68] = 8'h00;
mem[16'h2E69] = 8'h00;
mem[16'h2E6A] = 8'h00;
mem[16'h2E6B] = 8'h00;
mem[16'h2E6C] = 8'h00;
mem[16'h2E6D] = 8'h00;
mem[16'h2E6E] = 8'h00;
mem[16'h2E6F] = 8'h00;
mem[16'h2E70] = 8'h0F;
mem[16'h2E71] = 8'h40;
mem[16'h2E72] = 8'h07;
mem[16'h2E73] = 8'h00;
mem[16'h2E74] = 8'h00;
mem[16'h2E75] = 8'h00;
mem[16'h2E76] = 8'h00;
mem[16'h2E77] = 8'h2A;
mem[16'h2E78] = 8'h00;
mem[16'h2E79] = 8'h00;
mem[16'h2E7A] = 8'h00;
mem[16'h2E7B] = 8'h00;
mem[16'h2E7C] = 8'h00;
mem[16'h2E7D] = 8'h00;
mem[16'h2E7E] = 8'h00;
mem[16'h2E7F] = 8'h00;
mem[16'h2E80] = 8'hFD;
mem[16'h2E81] = 8'hD4;
mem[16'h2E82] = 8'hD2;
mem[16'h2E83] = 8'hCF;
mem[16'h2E84] = 8'hAA;
mem[16'h2E85] = 8'hAA;
mem[16'h2E86] = 8'hD5;
mem[16'h2E87] = 8'hAA;
mem[16'h2E88] = 8'hF5;
mem[16'h2E89] = 8'hD3;
mem[16'h2E8A] = 8'hCA;
mem[16'h2E8B] = 8'hBE;
mem[16'h2E8C] = 8'hAA;
mem[16'h2E8D] = 8'hA9;
mem[16'h2E8E] = 8'hD5;
mem[16'h2E8F] = 8'hAA;
mem[16'h2E90] = 8'hD5;
mem[16'h2E91] = 8'hCF;
mem[16'h2E92] = 8'hAA;
mem[16'h2E93] = 8'hFA;
mem[16'h2E94] = 8'hA9;
mem[16'h2E95] = 8'hA5;
mem[16'h2E96] = 8'hD5;
mem[16'h2E97] = 8'hAA;
mem[16'h2E98] = 8'hD5;
mem[16'h2E99] = 8'hBE;
mem[16'h2E9A] = 8'hAA;
mem[16'h2E9B] = 8'hE9;
mem[16'h2E9C] = 8'hA7;
mem[16'h2E9D] = 8'h95;
mem[16'h2E9E] = 8'hD5;
mem[16'h2E9F] = 8'hAA;
mem[16'h2EA0] = 8'hD5;
mem[16'h2EA1] = 8'hAA;
mem[16'h2EA2] = 8'hD5;
mem[16'h2EA3] = 8'hAA;
mem[16'h2EA4] = 8'h85;
mem[16'h2EA5] = 8'h00;
mem[16'h2EA6] = 8'h00;
mem[16'h2EA7] = 8'h00;
mem[16'h2EA8] = 8'h00;
mem[16'h2EA9] = 8'h00;
mem[16'h2EAA] = 8'h00;
mem[16'h2EAB] = 8'h00;
mem[16'h2EAC] = 8'h00;
mem[16'h2EAD] = 8'h00;
mem[16'h2EAE] = 8'h00;
mem[16'h2EAF] = 8'h00;
mem[16'h2EB0] = 8'h00;
mem[16'h2EB1] = 8'h00;
mem[16'h2EB2] = 8'h00;
mem[16'h2EB3] = 8'h00;
mem[16'h2EB4] = 8'h00;
mem[16'h2EB5] = 8'h00;
mem[16'h2EB6] = 8'h00;
mem[16'h2EB7] = 8'h00;
mem[16'h2EB8] = 8'h00;
mem[16'h2EB9] = 8'h00;
mem[16'h2EBA] = 8'h00;
mem[16'h2EBB] = 8'h00;
mem[16'h2EBC] = 8'h00;
mem[16'h2EBD] = 8'h00;
mem[16'h2EBE] = 8'h00;
mem[16'h2EBF] = 8'h00;
mem[16'h2EC0] = 8'h00;
mem[16'h2EC1] = 8'h00;
mem[16'h2EC2] = 8'h00;
mem[16'h2EC3] = 8'h00;
mem[16'h2EC4] = 8'h00;
mem[16'h2EC5] = 8'h00;
mem[16'h2EC6] = 8'h00;
mem[16'h2EC7] = 8'h00;
mem[16'h2EC8] = 8'h00;
mem[16'h2EC9] = 8'h00;
mem[16'h2ECA] = 8'h00;
mem[16'h2ECB] = 8'h00;
mem[16'h2ECC] = 8'h00;
mem[16'h2ECD] = 8'h00;
mem[16'h2ECE] = 8'h00;
mem[16'h2ECF] = 8'h2A;
mem[16'h2ED0] = 8'h00;
mem[16'h2ED1] = 8'h00;
mem[16'h2ED2] = 8'h00;
mem[16'h2ED3] = 8'h00;
mem[16'h2ED4] = 8'h0F;
mem[16'h2ED5] = 8'h40;
mem[16'h2ED6] = 8'h07;
mem[16'h2ED7] = 8'h00;
mem[16'h2ED8] = 8'h00;
mem[16'h2ED9] = 8'h00;
mem[16'h2EDA] = 8'h00;
mem[16'h2EDB] = 8'h00;
mem[16'h2EDC] = 8'h00;
mem[16'h2EDD] = 8'h00;
mem[16'h2EDE] = 8'h00;
mem[16'h2EDF] = 8'h00;
mem[16'h2EE0] = 8'h00;
mem[16'h2EE1] = 8'h00;
mem[16'h2EE2] = 8'h0F;
mem[16'h2EE3] = 8'h40;
mem[16'h2EE4] = 8'h07;
mem[16'h2EE5] = 8'h00;
mem[16'h2EE6] = 8'h00;
mem[16'h2EE7] = 8'h00;
mem[16'h2EE8] = 8'h00;
mem[16'h2EE9] = 8'h00;
mem[16'h2EEA] = 8'h00;
mem[16'h2EEB] = 8'h00;
mem[16'h2EEC] = 8'h00;
mem[16'h2EED] = 8'h00;
mem[16'h2EEE] = 8'h00;
mem[16'h2EEF] = 8'h00;
mem[16'h2EF0] = 8'h0F;
mem[16'h2EF1] = 8'h40;
mem[16'h2EF2] = 8'h07;
mem[16'h2EF3] = 8'h00;
mem[16'h2EF4] = 8'h00;
mem[16'h2EF5] = 8'h00;
mem[16'h2EF6] = 8'h00;
mem[16'h2EF7] = 8'h2A;
mem[16'h2EF8] = 8'h00;
mem[16'h2EF9] = 8'h00;
mem[16'h2EFA] = 8'h00;
mem[16'h2EFB] = 8'h00;
mem[16'h2EFC] = 8'h00;
mem[16'h2EFD] = 8'h00;
mem[16'h2EFE] = 8'h00;
mem[16'h2EFF] = 8'h00;
mem[16'h2F00] = 8'hEB;
mem[16'h2F01] = 8'hAA;
mem[16'h2F02] = 8'hD5;
mem[16'h2F03] = 8'hAA;
mem[16'h2F04] = 8'hD5;
mem[16'h2F05] = 8'hAA;
mem[16'h2F06] = 8'hD5;
mem[16'h2F07] = 8'hAA;
mem[16'h2F08] = 8'hD5;
mem[16'h2F09] = 8'hAA;
mem[16'h2F0A] = 8'hD5;
mem[16'h2F0B] = 8'hDA;
mem[16'h2F0C] = 8'hAA;
mem[16'h2F0D] = 8'hD5;
mem[16'h2F0E] = 8'hAA;
mem[16'h2F0F] = 8'hD5;
mem[16'h2F10] = 8'hAA;
mem[16'h2F11] = 8'hD5;
mem[16'h2F12] = 8'hAA;
mem[16'h2F13] = 8'hD5;
mem[16'h2F14] = 8'hAA;
mem[16'h2F15] = 8'hD5;
mem[16'h2F16] = 8'hAA;
mem[16'h2F17] = 8'hD5;
mem[16'h2F18] = 8'hAA;
mem[16'h2F19] = 8'hAD;
mem[16'h2F1A] = 8'hD5;
mem[16'h2F1B] = 8'hAA;
mem[16'h2F1C] = 8'hD5;
mem[16'h2F1D] = 8'hAA;
mem[16'h2F1E] = 8'hD5;
mem[16'h2F1F] = 8'hAA;
mem[16'h2F20] = 8'hD5;
mem[16'h2F21] = 8'hAA;
mem[16'h2F22] = 8'hD5;
mem[16'h2F23] = 8'hAA;
mem[16'h2F24] = 8'h85;
mem[16'h2F25] = 8'h00;
mem[16'h2F26] = 8'h74;
mem[16'h2F27] = 8'h17;
mem[16'h2F28] = 8'h00;
mem[16'h2F29] = 8'h00;
mem[16'h2F2A] = 8'h00;
mem[16'h2F2B] = 8'h03;
mem[16'h2F2C] = 8'h0C;
mem[16'h2F2D] = 8'h00;
mem[16'h2F2E] = 8'h00;
mem[16'h2F2F] = 8'h00;
mem[16'h2F30] = 8'h00;
mem[16'h2F31] = 8'h00;
mem[16'h2F32] = 8'h00;
mem[16'h2F33] = 8'h00;
mem[16'h2F34] = 8'h00;
mem[16'h2F35] = 8'h00;
mem[16'h2F36] = 8'h00;
mem[16'h2F37] = 8'h00;
mem[16'h2F38] = 8'h00;
mem[16'h2F39] = 8'h03;
mem[16'h2F3A] = 8'h0C;
mem[16'h2F3B] = 8'h00;
mem[16'h2F3C] = 8'h00;
mem[16'h2F3D] = 8'h00;
mem[16'h2F3E] = 8'h00;
mem[16'h2F3F] = 8'h00;
mem[16'h2F40] = 8'h00;
mem[16'h2F41] = 8'h00;
mem[16'h2F42] = 8'h00;
mem[16'h2F43] = 8'h00;
mem[16'h2F44] = 8'h00;
mem[16'h2F45] = 8'h00;
mem[16'h2F46] = 8'h00;
mem[16'h2F47] = 8'h00;
mem[16'h2F48] = 8'h00;
mem[16'h2F49] = 8'h00;
mem[16'h2F4A] = 8'h00;
mem[16'h2F4B] = 8'h00;
mem[16'h2F4C] = 8'h00;
mem[16'h2F4D] = 8'h00;
mem[16'h2F4E] = 8'h00;
mem[16'h2F4F] = 8'h2A;
mem[16'h2F50] = 8'h0A;
mem[16'h2F51] = 8'h04;
mem[16'h2F52] = 8'h2A;
mem[16'h2F53] = 8'h51;
mem[16'h2F54] = 8'h2A;
mem[16'h2F55] = 8'h54;
mem[16'h2F56] = 8'h22;
mem[16'h2F57] = 8'h54;
mem[16'h2F58] = 8'h0A;
mem[16'h2F59] = 8'h04;
mem[16'h2F5A] = 8'h2A;
mem[16'h2F5B] = 8'h51;
mem[16'h2F5C] = 8'h2A;
mem[16'h2F5D] = 8'h54;
mem[16'h2F5E] = 8'h22;
mem[16'h2F5F] = 8'h54;
mem[16'h2F60] = 8'h0A;
mem[16'h2F61] = 8'h04;
mem[16'h2F62] = 8'h40;
mem[16'h2F63] = 8'h01;
mem[16'h2F64] = 8'h2A;
mem[16'h2F65] = 8'h54;
mem[16'h2F66] = 8'h22;
mem[16'h2F67] = 8'h54;
mem[16'h2F68] = 8'h0A;
mem[16'h2F69] = 8'h04;
mem[16'h2F6A] = 8'h2A;
mem[16'h2F6B] = 8'h51;
mem[16'h2F6C] = 8'h2A;
mem[16'h2F6D] = 8'h54;
mem[16'h2F6E] = 8'h22;
mem[16'h2F6F] = 8'h54;
mem[16'h2F70] = 8'h0A;
mem[16'h2F71] = 8'h04;
mem[16'h2F72] = 8'h2A;
mem[16'h2F73] = 8'h51;
mem[16'h2F74] = 8'h0A;
mem[16'h2F75] = 8'h00;
mem[16'h2F76] = 8'h00;
mem[16'h2F77] = 8'h2A;
mem[16'h2F78] = 8'h00;
mem[16'h2F79] = 8'h00;
mem[16'h2F7A] = 8'h00;
mem[16'h2F7B] = 8'h00;
mem[16'h2F7C] = 8'h00;
mem[16'h2F7D] = 8'h00;
mem[16'h2F7E] = 8'h00;
mem[16'h2F7F] = 8'h00;
mem[16'h2F80] = 8'hEB;
mem[16'h2F81] = 8'hAA;
mem[16'h2F82] = 8'hD5;
mem[16'h2F83] = 8'hAA;
mem[16'h2F84] = 8'hD5;
mem[16'h2F85] = 8'hAA;
mem[16'h2F86] = 8'hD5;
mem[16'h2F87] = 8'hAA;
mem[16'h2F88] = 8'hD5;
mem[16'h2F89] = 8'hAA;
mem[16'h2F8A] = 8'hD5;
mem[16'h2F8B] = 8'hDA;
mem[16'h2F8C] = 8'hAA;
mem[16'h2F8D] = 8'hD5;
mem[16'h2F8E] = 8'hAA;
mem[16'h2F8F] = 8'hD5;
mem[16'h2F90] = 8'hAA;
mem[16'h2F91] = 8'hD5;
mem[16'h2F92] = 8'hAA;
mem[16'h2F93] = 8'hD5;
mem[16'h2F94] = 8'hAA;
mem[16'h2F95] = 8'hD5;
mem[16'h2F96] = 8'hAA;
mem[16'h2F97] = 8'hD5;
mem[16'h2F98] = 8'hAA;
mem[16'h2F99] = 8'hAD;
mem[16'h2F9A] = 8'hD5;
mem[16'h2F9B] = 8'hAA;
mem[16'h2F9C] = 8'hD5;
mem[16'h2F9D] = 8'hAA;
mem[16'h2F9E] = 8'hD5;
mem[16'h2F9F] = 8'hAA;
mem[16'h2FA0] = 8'hD5;
mem[16'h2FA1] = 8'hAA;
mem[16'h2FA2] = 8'hD5;
mem[16'h2FA3] = 8'hAA;
mem[16'h2FA4] = 8'h85;
mem[16'h2FA5] = 8'h00;
mem[16'h2FA6] = 8'h00;
mem[16'h2FA7] = 8'h00;
mem[16'h2FA8] = 8'h00;
mem[16'h2FA9] = 8'hF0;
mem[16'h2FAA] = 8'hC0;
mem[16'h2FAB] = 8'h83;
mem[16'h2FAC] = 8'h00;
mem[16'h2FAD] = 8'h00;
mem[16'h2FAE] = 8'h00;
mem[16'h2FAF] = 8'h00;
mem[16'h2FB0] = 8'h00;
mem[16'h2FB1] = 8'h00;
mem[16'h2FB2] = 8'h00;
mem[16'h2FB3] = 8'h00;
mem[16'h2FB4] = 8'h00;
mem[16'h2FB5] = 8'h00;
mem[16'h2FB6] = 8'h00;
mem[16'h2FB7] = 8'h00;
mem[16'h2FB8] = 8'h00;
mem[16'h2FB9] = 8'h00;
mem[16'h2FBA] = 8'h00;
mem[16'h2FBB] = 8'h00;
mem[16'h2FBC] = 8'h00;
mem[16'h2FBD] = 8'h00;
mem[16'h2FBE] = 8'h00;
mem[16'h2FBF] = 8'h00;
mem[16'h2FC0] = 8'h00;
mem[16'h2FC1] = 8'h00;
mem[16'h2FC2] = 8'h00;
mem[16'h2FC3] = 8'h00;
mem[16'h2FC4] = 8'h00;
mem[16'h2FC5] = 8'h00;
mem[16'h2FC6] = 8'h00;
mem[16'h2FC7] = 8'h00;
mem[16'h2FC8] = 8'h00;
mem[16'h2FC9] = 8'h00;
mem[16'h2FCA] = 8'h00;
mem[16'h2FCB] = 8'h00;
mem[16'h2FCC] = 8'h00;
mem[16'h2FCD] = 8'h00;
mem[16'h2FCE] = 8'h00;
mem[16'h2FCF] = 8'h2A;
mem[16'h2FD0] = 8'h0A;
mem[16'h2FD1] = 8'h04;
mem[16'h2FD2] = 8'h2A;
mem[16'h2FD3] = 8'h51;
mem[16'h2FD4] = 8'h2A;
mem[16'h2FD5] = 8'h54;
mem[16'h2FD6] = 8'h22;
mem[16'h2FD7] = 8'h54;
mem[16'h2FD8] = 8'h0A;
mem[16'h2FD9] = 8'h04;
mem[16'h2FDA] = 8'h2A;
mem[16'h2FDB] = 8'h51;
mem[16'h2FDC] = 8'h2A;
mem[16'h2FDD] = 8'h54;
mem[16'h2FDE] = 8'h22;
mem[16'h2FDF] = 8'h54;
mem[16'h2FE0] = 8'h0A;
mem[16'h2FE1] = 8'h04;
mem[16'h2FE2] = 8'h0E;
mem[16'h2FE3] = 8'h38;
mem[16'h2FE4] = 8'h2A;
mem[16'h2FE5] = 8'h54;
mem[16'h2FE6] = 8'h22;
mem[16'h2FE7] = 8'h54;
mem[16'h2FE8] = 8'h0A;
mem[16'h2FE9] = 8'h04;
mem[16'h2FEA] = 8'h2A;
mem[16'h2FEB] = 8'h51;
mem[16'h2FEC] = 8'h2A;
mem[16'h2FED] = 8'h54;
mem[16'h2FEE] = 8'h22;
mem[16'h2FEF] = 8'h54;
mem[16'h2FF0] = 8'h0A;
mem[16'h2FF1] = 8'h04;
mem[16'h2FF2] = 8'h2A;
mem[16'h2FF3] = 8'h51;
mem[16'h2FF4] = 8'h0A;
mem[16'h2FF5] = 8'h52;
mem[16'h2FF6] = 8'h00;
mem[16'h2FF7] = 8'h2A;
mem[16'h2FF8] = 8'h00;
mem[16'h2FF9] = 8'h00;
mem[16'h2FFA] = 8'h00;
mem[16'h2FFB] = 8'h00;
mem[16'h2FFC] = 8'h00;
mem[16'h2FFD] = 8'h00;
mem[16'h2FFE] = 8'h00;
mem[16'h2FFF] = 8'h00;
mem[16'h3000] = 8'h00;
mem[16'h3001] = 8'h42;
mem[16'h3002] = 8'h10;
mem[16'h3003] = 8'h00;
mem[16'h3004] = 8'h40;
mem[16'h3005] = 8'h02;
mem[16'h3006] = 8'h44;
mem[16'h3007] = 8'h02;
mem[16'h3008] = 8'h7E;
mem[16'h3009] = 8'h00;
mem[16'h300A] = 8'h42;
mem[16'h300B] = 8'h42;
mem[16'h300C] = 8'h42;
mem[16'h300D] = 8'h42;
mem[16'h300E] = 8'h42;
mem[16'h300F] = 8'h42;
mem[16'h3010] = 8'h00;
mem[16'h3011] = 8'h00;
mem[16'h3012] = 8'h00;
mem[16'h3013] = 8'h00;
mem[16'h3014] = 8'h10;
mem[16'h3015] = 8'h44;
mem[16'h3016] = 8'h42;
mem[16'h3017] = 8'h02;
mem[16'h3018] = 8'h00;
mem[16'h3019] = 8'h40;
mem[16'h301A] = 8'h02;
mem[16'h301B] = 8'h44;
mem[16'h301C] = 8'h02;
mem[16'h301D] = 8'h7E;
mem[16'h301E] = 8'h00;
mem[16'h301F] = 8'h42;
mem[16'h3020] = 8'h42;
mem[16'h3021] = 8'h42;
mem[16'h3022] = 8'h42;
mem[16'h3023] = 8'h42;
mem[16'h3024] = 8'h42;
mem[16'h3025] = 8'h00;
mem[16'h3026] = 8'h60;
mem[16'h3027] = 8'h03;
mem[16'h3028] = 8'hD5;
mem[16'h3029] = 8'hAA;
mem[16'h302A] = 8'hD5;
mem[16'h302B] = 8'hAA;
mem[16'h302C] = 8'hB5;
mem[16'h302D] = 8'hD5;
mem[16'h302E] = 8'hAA;
mem[16'h302F] = 8'hD5;
mem[16'h3030] = 8'hAA;
mem[16'h3031] = 8'hD5;
mem[16'h3032] = 8'hAA;
mem[16'h3033] = 8'hD5;
mem[16'h3034] = 8'hD6;
mem[16'h3035] = 8'hAA;
mem[16'h3036] = 8'hD5;
mem[16'h3037] = 8'hAA;
mem[16'h3038] = 8'hD5;
mem[16'h3039] = 8'hD5;
mem[16'h303A] = 8'hAA;
mem[16'h303B] = 8'hD5;
mem[16'h303C] = 8'hAA;
mem[16'h303D] = 8'hD5;
mem[16'h303E] = 8'hAA;
mem[16'h303F] = 8'hD5;
mem[16'h3040] = 8'hDA;
mem[16'h3041] = 8'hAA;
mem[16'h3042] = 8'hD5;
mem[16'h3043] = 8'hAA;
mem[16'h3044] = 8'hAB;
mem[16'h3045] = 8'hD5;
mem[16'h3046] = 8'hAA;
mem[16'h3047] = 8'hD5;
mem[16'h3048] = 8'hAA;
mem[16'h3049] = 8'hD5;
mem[16'h304A] = 8'hAA;
mem[16'h304B] = 8'hB5;
mem[16'h304C] = 8'h85;
mem[16'h304D] = 8'h00;
mem[16'h304E] = 8'h00;
mem[16'h304F] = 8'h00;
mem[16'h3050] = 8'h00;
mem[16'h3051] = 8'h00;
mem[16'h3052] = 8'h00;
mem[16'h3053] = 8'h00;
mem[16'h3054] = 8'h00;
mem[16'h3055] = 8'h00;
mem[16'h3056] = 8'h00;
mem[16'h3057] = 8'h00;
mem[16'h3058] = 8'h00;
mem[16'h3059] = 8'h00;
mem[16'h305A] = 8'h00;
mem[16'h305B] = 8'h00;
mem[16'h305C] = 8'h00;
mem[16'h305D] = 8'h00;
mem[16'h305E] = 8'h00;
mem[16'h305F] = 8'h00;
mem[16'h3060] = 8'h00;
mem[16'h3061] = 8'h00;
mem[16'h3062] = 8'h00;
mem[16'h3063] = 8'h00;
mem[16'h3064] = 8'h00;
mem[16'h3065] = 8'h00;
mem[16'h3066] = 8'h00;
mem[16'h3067] = 8'h00;
mem[16'h3068] = 8'h00;
mem[16'h3069] = 8'h00;
mem[16'h306A] = 8'h00;
mem[16'h306B] = 8'h00;
mem[16'h306C] = 8'h00;
mem[16'h306D] = 8'h00;
mem[16'h306E] = 8'h00;
mem[16'h306F] = 8'h00;
mem[16'h3070] = 8'h00;
mem[16'h3071] = 8'h00;
mem[16'h3072] = 8'h00;
mem[16'h3073] = 8'h00;
mem[16'h3074] = 8'h00;
mem[16'h3075] = 8'h00;
mem[16'h3076] = 8'h00;
mem[16'h3077] = 8'h2A;
mem[16'h3078] = 8'h00;
mem[16'h3079] = 8'h00;
mem[16'h307A] = 8'h00;
mem[16'h307B] = 8'h00;
mem[16'h307C] = 8'h00;
mem[16'h307D] = 8'h00;
mem[16'h307E] = 8'h00;
mem[16'h307F] = 8'h00;
mem[16'h3080] = 8'h2A;
mem[16'h3081] = 8'h45;
mem[16'h3082] = 8'h2A;
mem[16'h3083] = 8'hAA;
mem[16'h3084] = 8'hD5;
mem[16'h3085] = 8'h41;
mem[16'h3086] = 8'h20;
mem[16'h3087] = 8'h15;
mem[16'h3088] = 8'h2A;
mem[16'h3089] = 8'h45;
mem[16'h308A] = 8'hD5;
mem[16'h308B] = 8'hAA;
mem[16'h308C] = 8'h2A;
mem[16'h308D] = 8'h41;
mem[16'h308E] = 8'h20;
mem[16'h308F] = 8'h15;
mem[16'h3090] = 8'hD5;
mem[16'h3091] = 8'hAA;
mem[16'h3092] = 8'h2A;
mem[16'h3093] = 8'h44;
mem[16'h3094] = 8'h2A;
mem[16'h3095] = 8'h41;
mem[16'h3096] = 8'h20;
mem[16'h3097] = 8'hAA;
mem[16'h3098] = 8'hD5;
mem[16'h3099] = 8'h45;
mem[16'h309A] = 8'h2A;
mem[16'h309B] = 8'h44;
mem[16'h309C] = 8'h2A;
mem[16'h309D] = 8'hAA;
mem[16'h309E] = 8'hD5;
mem[16'h309F] = 8'h15;
mem[16'h30A0] = 8'h2A;
mem[16'h30A1] = 8'h45;
mem[16'h30A2] = 8'h2A;
mem[16'h30A3] = 8'h44;
mem[16'h30A4] = 8'h0A;
mem[16'h30A5] = 8'h00;
mem[16'h30A6] = 8'h44;
mem[16'h30A7] = 8'h12;
mem[16'h30A8] = 8'hD5;
mem[16'h30A9] = 8'hAA;
mem[16'h30AA] = 8'hD5;
mem[16'h30AB] = 8'hAA;
mem[16'h30AC] = 8'hD5;
mem[16'h30AD] = 8'h8A;
mem[16'h30AE] = 8'hD5;
mem[16'h30AF] = 8'hAA;
mem[16'h30B0] = 8'hD1;
mem[16'h30B1] = 8'hAA;
mem[16'h30B2] = 8'h95;
mem[16'h30B3] = 8'hAA;
mem[16'h30B4] = 8'hD5;
mem[16'h30B5] = 8'hAA;
mem[16'h30B6] = 8'hD5;
mem[16'h30B7] = 8'hAA;
mem[16'h30B8] = 8'hD5;
mem[16'h30B9] = 8'hAA;
mem[16'h30BA] = 8'hD5;
mem[16'h30BB] = 8'hAA;
mem[16'h30BC] = 8'hC5;
mem[16'h30BD] = 8'hAA;
mem[16'h30BE] = 8'hD5;
mem[16'h30BF] = 8'hA8;
mem[16'h30C0] = 8'hD5;
mem[16'h30C1] = 8'h8A;
mem[16'h30C2] = 8'hD5;
mem[16'h30C3] = 8'hAA;
mem[16'h30C4] = 8'hD5;
mem[16'h30C5] = 8'hAA;
mem[16'h30C6] = 8'hD5;
mem[16'h30C7] = 8'hAA;
mem[16'h30C8] = 8'hD5;
mem[16'h30C9] = 8'hAA;
mem[16'h30CA] = 8'hD5;
mem[16'h30CB] = 8'hAA;
mem[16'h30CC] = 8'h85;
mem[16'h30CD] = 8'h00;
mem[16'h30CE] = 8'h00;
mem[16'h30CF] = 8'h2A;
mem[16'h30D0] = 8'h00;
mem[16'h30D1] = 8'h00;
mem[16'h30D2] = 8'h00;
mem[16'h30D3] = 8'h00;
mem[16'h30D4] = 8'h00;
mem[16'h30D5] = 8'h56;
mem[16'h30D6] = 8'h2A;
mem[16'h30D7] = 8'h0F;
mem[16'h30D8] = 8'h00;
mem[16'h30D9] = 8'h00;
mem[16'h30DA] = 8'h00;
mem[16'h30DB] = 8'h00;
mem[16'h30DC] = 8'h00;
mem[16'h30DD] = 8'h00;
mem[16'h30DE] = 8'h00;
mem[16'h30DF] = 8'h00;
mem[16'h30E0] = 8'h00;
mem[16'h30E1] = 8'h56;
mem[16'h30E2] = 8'h2A;
mem[16'h30E3] = 8'h0F;
mem[16'h30E4] = 8'h00;
mem[16'h30E5] = 8'h00;
mem[16'h30E6] = 8'h00;
mem[16'h30E7] = 8'h00;
mem[16'h30E8] = 8'h00;
mem[16'h30E9] = 8'h00;
mem[16'h30EA] = 8'h00;
mem[16'h30EB] = 8'h00;
mem[16'h30EC] = 8'h00;
mem[16'h30ED] = 8'h56;
mem[16'h30EE] = 8'h2A;
mem[16'h30EF] = 8'h0F;
mem[16'h30F0] = 8'h00;
mem[16'h30F1] = 8'h00;
mem[16'h30F2] = 8'h00;
mem[16'h30F3] = 8'h00;
mem[16'h30F4] = 8'h00;
mem[16'h30F5] = 8'h00;
mem[16'h30F6] = 8'h00;
mem[16'h30F7] = 8'h2A;
mem[16'h30F8] = 8'h00;
mem[16'h30F9] = 8'h00;
mem[16'h30FA] = 8'h00;
mem[16'h30FB] = 8'h00;
mem[16'h30FC] = 8'h00;
mem[16'h30FD] = 8'h00;
mem[16'h30FE] = 8'h00;
mem[16'h30FF] = 8'h00;
mem[16'h3100] = 8'hD5;
mem[16'h3101] = 8'hAA;
mem[16'h3102] = 8'hD5;
mem[16'h3103] = 8'hAA;
mem[16'h3104] = 8'hD5;
mem[16'h3105] = 8'hAA;
mem[16'h3106] = 8'hD5;
mem[16'h3107] = 8'hAA;
mem[16'h3108] = 8'hD5;
mem[16'h3109] = 8'hAA;
mem[16'h310A] = 8'hD5;
mem[16'h310B] = 8'hAA;
mem[16'h310C] = 8'hD5;
mem[16'h310D] = 8'hAA;
mem[16'h310E] = 8'hD5;
mem[16'h310F] = 8'hAA;
mem[16'h3110] = 8'hD5;
mem[16'h3111] = 8'hAA;
mem[16'h3112] = 8'hD5;
mem[16'h3113] = 8'hAA;
mem[16'h3114] = 8'hD5;
mem[16'h3115] = 8'hAA;
mem[16'h3116] = 8'hD5;
mem[16'h3117] = 8'hAA;
mem[16'h3118] = 8'hD5;
mem[16'h3119] = 8'hAA;
mem[16'h311A] = 8'hD5;
mem[16'h311B] = 8'hAA;
mem[16'h311C] = 8'hD5;
mem[16'h311D] = 8'hAA;
mem[16'h311E] = 8'hD5;
mem[16'h311F] = 8'hAA;
mem[16'h3120] = 8'hD5;
mem[16'h3121] = 8'hAA;
mem[16'h3122] = 8'hD5;
mem[16'h3123] = 8'hAA;
mem[16'h3124] = 8'h85;
mem[16'h3125] = 8'h00;
mem[16'h3126] = 8'h40;
mem[16'h3127] = 8'h01;
mem[16'h3128] = 8'hD5;
mem[16'h3129] = 8'hAA;
mem[16'h312A] = 8'hD5;
mem[16'h312B] = 8'hAA;
mem[16'h312C] = 8'hD5;
mem[16'h312D] = 8'hCA;
mem[16'h312E] = 8'hC2;
mem[16'h312F] = 8'hAA;
mem[16'h3130] = 8'hA9;
mem[16'h3131] = 8'hA8;
mem[16'h3132] = 8'h95;
mem[16'h3133] = 8'h85;
mem[16'h3134] = 8'hD5;
mem[16'h3135] = 8'hAA;
mem[16'h3136] = 8'hD5;
mem[16'h3137] = 8'hAA;
mem[16'h3138] = 8'hD5;
mem[16'h3139] = 8'hAA;
mem[16'h313A] = 8'hD5;
mem[16'h313B] = 8'hAA;
mem[16'h313C] = 8'hA5;
mem[16'h313D] = 8'hA1;
mem[16'h313E] = 8'hD5;
mem[16'h313F] = 8'h94;
mem[16'h3140] = 8'hD4;
mem[16'h3141] = 8'hCA;
mem[16'h3142] = 8'hC2;
mem[16'h3143] = 8'hAA;
mem[16'h3144] = 8'hD5;
mem[16'h3145] = 8'hAA;
mem[16'h3146] = 8'hD5;
mem[16'h3147] = 8'hAA;
mem[16'h3148] = 8'hD5;
mem[16'h3149] = 8'hAA;
mem[16'h314A] = 8'hD5;
mem[16'h314B] = 8'hAA;
mem[16'h314C] = 8'h85;
mem[16'h314D] = 8'h00;
mem[16'h314E] = 8'h00;
mem[16'h314F] = 8'h2A;
mem[16'h3150] = 8'h00;
mem[16'h3151] = 8'h00;
mem[16'h3152] = 8'h00;
mem[16'h3153] = 8'h00;
mem[16'h3154] = 8'h00;
mem[16'h3155] = 8'h00;
mem[16'h3156] = 8'h00;
mem[16'h3157] = 8'h00;
mem[16'h3158] = 8'h00;
mem[16'h3159] = 8'h00;
mem[16'h315A] = 8'h00;
mem[16'h315B] = 8'h00;
mem[16'h315C] = 8'h00;
mem[16'h315D] = 8'h00;
mem[16'h315E] = 8'h00;
mem[16'h315F] = 8'h00;
mem[16'h3160] = 8'h00;
mem[16'h3161] = 8'h00;
mem[16'h3162] = 8'h00;
mem[16'h3163] = 8'h00;
mem[16'h3164] = 8'h00;
mem[16'h3165] = 8'h00;
mem[16'h3166] = 8'h00;
mem[16'h3167] = 8'h00;
mem[16'h3168] = 8'h00;
mem[16'h3169] = 8'h00;
mem[16'h316A] = 8'h00;
mem[16'h316B] = 8'h00;
mem[16'h316C] = 8'h00;
mem[16'h316D] = 8'h00;
mem[16'h316E] = 8'h00;
mem[16'h316F] = 8'h00;
mem[16'h3170] = 8'h00;
mem[16'h3171] = 8'h00;
mem[16'h3172] = 8'h00;
mem[16'h3173] = 8'h00;
mem[16'h3174] = 8'h00;
mem[16'h3175] = 8'h00;
mem[16'h3176] = 8'h00;
mem[16'h3177] = 8'h2A;
mem[16'h3178] = 8'h00;
mem[16'h3179] = 8'h00;
mem[16'h317A] = 8'h00;
mem[16'h317B] = 8'h00;
mem[16'h317C] = 8'h00;
mem[16'h317D] = 8'h00;
mem[16'h317E] = 8'h00;
mem[16'h317F] = 8'h00;
mem[16'h3180] = 8'hD5;
mem[16'h3181] = 8'hAA;
mem[16'h3182] = 8'hD5;
mem[16'h3183] = 8'hAA;
mem[16'h3184] = 8'hD5;
mem[16'h3185] = 8'hAA;
mem[16'h3186] = 8'hAB;
mem[16'h3187] = 8'hD5;
mem[16'h3188] = 8'hAA;
mem[16'h3189] = 8'hD5;
mem[16'h318A] = 8'hAA;
mem[16'h318B] = 8'hD5;
mem[16'h318C] = 8'hAA;
mem[16'h318D] = 8'hD5;
mem[16'h318E] = 8'hAA;
mem[16'h318F] = 8'hD5;
mem[16'h3190] = 8'hD5;
mem[16'h3191] = 8'hAA;
mem[16'h3192] = 8'hAD;
mem[16'h3193] = 8'hD5;
mem[16'h3194] = 8'hAA;
mem[16'h3195] = 8'hD5;
mem[16'h3196] = 8'hAA;
mem[16'h3197] = 8'hD5;
mem[16'h3198] = 8'hAA;
mem[16'h3199] = 8'hD5;
mem[16'h319A] = 8'hAA;
mem[16'h319B] = 8'hD5;
mem[16'h319C] = 8'hD6;
mem[16'h319D] = 8'hAA;
mem[16'h319E] = 8'hD5;
mem[16'h319F] = 8'hAA;
mem[16'h31A0] = 8'hD5;
mem[16'h31A1] = 8'hAA;
mem[16'h31A2] = 8'hD5;
mem[16'h31A3] = 8'hAA;
mem[16'h31A4] = 8'h85;
mem[16'h31A5] = 8'h00;
mem[16'h31A6] = 8'h0E;
mem[16'h31A7] = 8'h38;
mem[16'h31A8] = 8'h22;
mem[16'h31A9] = 8'h15;
mem[16'h31AA] = 8'h22;
mem[16'h31AB] = 8'h55;
mem[16'h31AC] = 8'h20;
mem[16'h31AD] = 8'h50;
mem[16'h31AE] = 8'h0A;
mem[16'h31AF] = 8'h55;
mem[16'h31B0] = 8'h22;
mem[16'h31B1] = 8'h15;
mem[16'h31B2] = 8'h22;
mem[16'h31B3] = 8'h55;
mem[16'h31B4] = 8'h20;
mem[16'h31B5] = 8'h50;
mem[16'h31B6] = 8'h0A;
mem[16'h31B7] = 8'h55;
mem[16'h31B8] = 8'h22;
mem[16'h31B9] = 8'h15;
mem[16'h31BA] = 8'h22;
mem[16'h31BB] = 8'h55;
mem[16'h31BC] = 8'h20;
mem[16'h31BD] = 8'h50;
mem[16'h31BE] = 8'h0A;
mem[16'h31BF] = 8'h55;
mem[16'h31C0] = 8'h22;
mem[16'h31C1] = 8'h15;
mem[16'h31C2] = 8'h22;
mem[16'h31C3] = 8'h55;
mem[16'h31C4] = 8'h20;
mem[16'h31C5] = 8'h50;
mem[16'h31C6] = 8'h0A;
mem[16'h31C7] = 8'h55;
mem[16'h31C8] = 8'h22;
mem[16'h31C9] = 8'h15;
mem[16'h31CA] = 8'h22;
mem[16'h31CB] = 8'h55;
mem[16'h31CC] = 8'h00;
mem[16'h31CD] = 8'h00;
mem[16'h31CE] = 8'h00;
mem[16'h31CF] = 8'h2A;
mem[16'h31D0] = 8'h00;
mem[16'h31D1] = 8'hD8;
mem[16'h31D2] = 8'h8D;
mem[16'h31D3] = 8'h82;
mem[16'h31D4] = 8'h00;
mem[16'h31D5] = 8'h00;
mem[16'h31D6] = 8'h00;
mem[16'h31D7] = 8'h00;
mem[16'h31D8] = 8'h00;
mem[16'h31D9] = 8'h00;
mem[16'h31DA] = 8'h00;
mem[16'h31DB] = 8'hC0;
mem[16'h31DC] = 8'hED;
mem[16'h31DD] = 8'h90;
mem[16'h31DE] = 8'h00;
mem[16'h31DF] = 8'h00;
mem[16'h31E0] = 8'h00;
mem[16'h31E1] = 8'h00;
mem[16'h31E2] = 8'h00;
mem[16'h31E3] = 8'h00;
mem[16'h31E4] = 8'h00;
mem[16'h31E5] = 8'h00;
mem[16'h31E6] = 8'hEC;
mem[16'h31E7] = 8'h86;
mem[16'h31E8] = 8'h81;
mem[16'h31E9] = 8'h00;
mem[16'h31EA] = 8'h00;
mem[16'h31EB] = 8'h00;
mem[16'h31EC] = 8'h00;
mem[16'h31ED] = 8'h00;
mem[16'h31EE] = 8'h00;
mem[16'h31EF] = 8'h00;
mem[16'h31F0] = 8'h00;
mem[16'h31F1] = 8'h00;
mem[16'h31F2] = 8'h00;
mem[16'h31F3] = 8'h00;
mem[16'h31F4] = 8'h00;
mem[16'h31F5] = 8'h00;
mem[16'h31F6] = 8'h00;
mem[16'h31F7] = 8'h2A;
mem[16'h31F8] = 8'h00;
mem[16'h31F9] = 8'h00;
mem[16'h31FA] = 8'h00;
mem[16'h31FB] = 8'h00;
mem[16'h31FC] = 8'h00;
mem[16'h31FD] = 8'h00;
mem[16'h31FE] = 8'h00;
mem[16'h31FF] = 8'h00;
mem[16'h3200] = 8'hD5;
mem[16'h3201] = 8'hAA;
mem[16'h3202] = 8'hD5;
mem[16'h3203] = 8'hAA;
mem[16'h3204] = 8'hD5;
mem[16'h3205] = 8'hAA;
mem[16'h3206] = 8'hD5;
mem[16'h3207] = 8'hAA;
mem[16'h3208] = 8'hD5;
mem[16'h3209] = 8'hAA;
mem[16'h320A] = 8'hD5;
mem[16'h320B] = 8'hAA;
mem[16'h320C] = 8'hD5;
mem[16'h320D] = 8'hAA;
mem[16'h320E] = 8'hD5;
mem[16'h320F] = 8'hAA;
mem[16'h3210] = 8'hD5;
mem[16'h3211] = 8'hAA;
mem[16'h3212] = 8'hD5;
mem[16'h3213] = 8'hAA;
mem[16'h3214] = 8'hD5;
mem[16'h3215] = 8'hAA;
mem[16'h3216] = 8'hD5;
mem[16'h3217] = 8'hAA;
mem[16'h3218] = 8'hD5;
mem[16'h3219] = 8'hAA;
mem[16'h321A] = 8'hD5;
mem[16'h321B] = 8'hAA;
mem[16'h321C] = 8'hD5;
mem[16'h321D] = 8'hAA;
mem[16'h321E] = 8'hD5;
mem[16'h321F] = 8'hAA;
mem[16'h3220] = 8'hD5;
mem[16'h3221] = 8'hAA;
mem[16'h3222] = 8'hD5;
mem[16'h3223] = 8'hAA;
mem[16'h3224] = 8'h85;
mem[16'h3225] = 8'h00;
mem[16'h3226] = 8'h70;
mem[16'h3227] = 8'h07;
mem[16'h3228] = 8'h22;
mem[16'h3229] = 8'h15;
mem[16'h322A] = 8'h22;
mem[16'h322B] = 8'h55;
mem[16'h322C] = 8'h20;
mem[16'h322D] = 8'h50;
mem[16'h322E] = 8'h0A;
mem[16'h322F] = 8'h55;
mem[16'h3230] = 8'h22;
mem[16'h3231] = 8'h15;
mem[16'h3232] = 8'h22;
mem[16'h3233] = 8'h55;
mem[16'h3234] = 8'h20;
mem[16'h3235] = 8'h50;
mem[16'h3236] = 8'h0A;
mem[16'h3237] = 8'h55;
mem[16'h3238] = 8'h22;
mem[16'h3239] = 8'h15;
mem[16'h323A] = 8'h22;
mem[16'h323B] = 8'h55;
mem[16'h323C] = 8'h20;
mem[16'h323D] = 8'h50;
mem[16'h323E] = 8'h0A;
mem[16'h323F] = 8'h55;
mem[16'h3240] = 8'h22;
mem[16'h3241] = 8'h15;
mem[16'h3242] = 8'h22;
mem[16'h3243] = 8'h55;
mem[16'h3244] = 8'h20;
mem[16'h3245] = 8'h50;
mem[16'h3246] = 8'h0A;
mem[16'h3247] = 8'h55;
mem[16'h3248] = 8'h22;
mem[16'h3249] = 8'h15;
mem[16'h324A] = 8'h22;
mem[16'h324B] = 8'h55;
mem[16'h324C] = 8'h00;
mem[16'h324D] = 8'h00;
mem[16'h324E] = 8'h00;
mem[16'h324F] = 8'h2A;
mem[16'h3250] = 8'h00;
mem[16'h3251] = 8'h00;
mem[16'h3252] = 8'h00;
mem[16'h3253] = 8'h00;
mem[16'h3254] = 8'h4F;
mem[16'h3255] = 8'h4A;
mem[16'h3256] = 8'h07;
mem[16'h3257] = 8'h00;
mem[16'h3258] = 8'h00;
mem[16'h3259] = 8'h00;
mem[16'h325A] = 8'h00;
mem[16'h325B] = 8'h00;
mem[16'h325C] = 8'h00;
mem[16'h325D] = 8'h00;
mem[16'h325E] = 8'h00;
mem[16'h325F] = 8'h00;
mem[16'h3260] = 8'h00;
mem[16'h3261] = 8'h00;
mem[16'h3262] = 8'h4F;
mem[16'h3263] = 8'h4A;
mem[16'h3264] = 8'h07;
mem[16'h3265] = 8'h00;
mem[16'h3266] = 8'h00;
mem[16'h3267] = 8'h00;
mem[16'h3268] = 8'h00;
mem[16'h3269] = 8'h00;
mem[16'h326A] = 8'h00;
mem[16'h326B] = 8'h00;
mem[16'h326C] = 8'h00;
mem[16'h326D] = 8'h00;
mem[16'h326E] = 8'h00;
mem[16'h326F] = 8'h00;
mem[16'h3270] = 8'h4F;
mem[16'h3271] = 8'h4A;
mem[16'h3272] = 8'h07;
mem[16'h3273] = 8'h00;
mem[16'h3274] = 8'h00;
mem[16'h3275] = 8'h00;
mem[16'h3276] = 8'h00;
mem[16'h3277] = 8'h2A;
mem[16'h3278] = 8'h00;
mem[16'h3279] = 8'h00;
mem[16'h327A] = 8'h00;
mem[16'h327B] = 8'h00;
mem[16'h327C] = 8'h00;
mem[16'h327D] = 8'h00;
mem[16'h327E] = 8'h00;
mem[16'h327F] = 8'h00;
mem[16'h3280] = 8'hB5;
mem[16'h3281] = 8'hD5;
mem[16'h3282] = 8'hD4;
mem[16'h3283] = 8'hD6;
mem[16'h3284] = 8'hCA;
mem[16'h3285] = 8'hAA;
mem[16'h3286] = 8'hD5;
mem[16'h3287] = 8'hAA;
mem[16'h3288] = 8'hD5;
mem[16'h3289] = 8'hD5;
mem[16'h328A] = 8'hD2;
mem[16'h328B] = 8'hDA;
mem[16'h328C] = 8'hAA;
mem[16'h328D] = 8'hAA;
mem[16'h328E] = 8'hD5;
mem[16'h328F] = 8'hAA;
mem[16'h3290] = 8'hD5;
mem[16'h3291] = 8'hD6;
mem[16'h3292] = 8'hCA;
mem[16'h3293] = 8'hEA;
mem[16'h3294] = 8'hAA;
mem[16'h3295] = 8'hA9;
mem[16'h3296] = 8'hD5;
mem[16'h3297] = 8'hAA;
mem[16'h3298] = 8'hD5;
mem[16'h3299] = 8'hDA;
mem[16'h329A] = 8'hAA;
mem[16'h329B] = 8'hAA;
mem[16'h329C] = 8'hAB;
mem[16'h329D] = 8'hA5;
mem[16'h329E] = 8'hD5;
mem[16'h329F] = 8'hAA;
mem[16'h32A0] = 8'hD5;
mem[16'h32A1] = 8'hAA;
mem[16'h32A2] = 8'hD5;
mem[16'h32A3] = 8'hAA;
mem[16'h32A4] = 8'h85;
mem[16'h32A5] = 8'h00;
mem[16'h32A6] = 8'h00;
mem[16'h32A7] = 8'h00;
mem[16'h32A8] = 8'h00;
mem[16'h32A9] = 8'h00;
mem[16'h32AA] = 8'h00;
mem[16'h32AB] = 8'h03;
mem[16'h32AC] = 8'h0C;
mem[16'h32AD] = 8'h00;
mem[16'h32AE] = 8'h00;
mem[16'h32AF] = 8'h00;
mem[16'h32B0] = 8'h00;
mem[16'h32B1] = 8'h00;
mem[16'h32B2] = 8'h00;
mem[16'h32B3] = 8'h00;
mem[16'h32B4] = 8'h00;
mem[16'h32B5] = 8'h00;
mem[16'h32B6] = 8'h00;
mem[16'h32B7] = 8'h00;
mem[16'h32B8] = 8'h00;
mem[16'h32B9] = 8'h03;
mem[16'h32BA] = 8'h0C;
mem[16'h32BB] = 8'h00;
mem[16'h32BC] = 8'h00;
mem[16'h32BD] = 8'h00;
mem[16'h32BE] = 8'h00;
mem[16'h32BF] = 8'h00;
mem[16'h32C0] = 8'h00;
mem[16'h32C1] = 8'h00;
mem[16'h32C2] = 8'h00;
mem[16'h32C3] = 8'h00;
mem[16'h32C4] = 8'h00;
mem[16'h32C5] = 8'h00;
mem[16'h32C6] = 8'h00;
mem[16'h32C7] = 8'h00;
mem[16'h32C8] = 8'h00;
mem[16'h32C9] = 8'h00;
mem[16'h32CA] = 8'h00;
mem[16'h32CB] = 8'h00;
mem[16'h32CC] = 8'h00;
mem[16'h32CD] = 8'h00;
mem[16'h32CE] = 8'h00;
mem[16'h32CF] = 8'h2A;
mem[16'h32D0] = 8'h00;
mem[16'h32D1] = 8'h00;
mem[16'h32D2] = 8'h00;
mem[16'h32D3] = 8'h00;
mem[16'h32D4] = 8'h00;
mem[16'h32D5] = 8'h00;
mem[16'h32D6] = 8'h00;
mem[16'h32D7] = 8'h00;
mem[16'h32D8] = 8'h00;
mem[16'h32D9] = 8'h00;
mem[16'h32DA] = 8'h00;
mem[16'h32DB] = 8'h00;
mem[16'h32DC] = 8'h00;
mem[16'h32DD] = 8'h00;
mem[16'h32DE] = 8'h00;
mem[16'h32DF] = 8'h00;
mem[16'h32E0] = 8'h00;
mem[16'h32E1] = 8'h00;
mem[16'h32E2] = 8'h00;
mem[16'h32E3] = 8'h00;
mem[16'h32E4] = 8'h00;
mem[16'h32E5] = 8'h00;
mem[16'h32E6] = 8'h00;
mem[16'h32E7] = 8'h00;
mem[16'h32E8] = 8'h00;
mem[16'h32E9] = 8'h00;
mem[16'h32EA] = 8'h00;
mem[16'h32EB] = 8'h00;
mem[16'h32EC] = 8'h00;
mem[16'h32ED] = 8'h00;
mem[16'h32EE] = 8'h00;
mem[16'h32EF] = 8'h00;
mem[16'h32F0] = 8'h00;
mem[16'h32F1] = 8'h00;
mem[16'h32F2] = 8'h00;
mem[16'h32F3] = 8'h00;
mem[16'h32F4] = 8'h00;
mem[16'h32F5] = 8'h00;
mem[16'h32F6] = 8'h00;
mem[16'h32F7] = 8'h2A;
mem[16'h32F8] = 8'h00;
mem[16'h32F9] = 8'h00;
mem[16'h32FA] = 8'h00;
mem[16'h32FB] = 8'h00;
mem[16'h32FC] = 8'h00;
mem[16'h32FD] = 8'h00;
mem[16'h32FE] = 8'h00;
mem[16'h32FF] = 8'h00;
mem[16'h3300] = 8'hAB;
mem[16'h3301] = 8'hAB;
mem[16'h3302] = 8'hD5;
mem[16'h3303] = 8'hAA;
mem[16'h3304] = 8'hD5;
mem[16'h3305] = 8'hAA;
mem[16'h3306] = 8'hD5;
mem[16'h3307] = 8'hAA;
mem[16'h3308] = 8'hD5;
mem[16'h3309] = 8'hAA;
mem[16'h330A] = 8'hD5;
mem[16'h330B] = 8'hD6;
mem[16'h330C] = 8'hAA;
mem[16'h330D] = 8'hD5;
mem[16'h330E] = 8'hAA;
mem[16'h330F] = 8'hD5;
mem[16'h3310] = 8'hAA;
mem[16'h3311] = 8'hD5;
mem[16'h3312] = 8'hAA;
mem[16'h3313] = 8'hD5;
mem[16'h3314] = 8'hAA;
mem[16'h3315] = 8'hD5;
mem[16'h3316] = 8'hAA;
mem[16'h3317] = 8'hD5;
mem[16'h3318] = 8'hAA;
mem[16'h3319] = 8'hB5;
mem[16'h331A] = 8'hD5;
mem[16'h331B] = 8'hAA;
mem[16'h331C] = 8'hD5;
mem[16'h331D] = 8'hAA;
mem[16'h331E] = 8'hD5;
mem[16'h331F] = 8'hAA;
mem[16'h3320] = 8'hD5;
mem[16'h3321] = 8'hAA;
mem[16'h3322] = 8'hD5;
mem[16'h3323] = 8'hAA;
mem[16'h3324] = 8'h85;
mem[16'h3325] = 8'h00;
mem[16'h3326] = 8'h7C;
mem[16'h3327] = 8'h1F;
mem[16'h3328] = 8'h00;
mem[16'h3329] = 8'h00;
mem[16'h332A] = 8'h00;
mem[16'h332B] = 8'h00;
mem[16'h332C] = 8'h00;
mem[16'h332D] = 8'h00;
mem[16'h332E] = 8'h00;
mem[16'h332F] = 8'h00;
mem[16'h3330] = 8'h00;
mem[16'h3331] = 8'h00;
mem[16'h3332] = 8'h00;
mem[16'h3333] = 8'h00;
mem[16'h3334] = 8'h00;
mem[16'h3335] = 8'h00;
mem[16'h3336] = 8'h00;
mem[16'h3337] = 8'h00;
mem[16'h3338] = 8'h00;
mem[16'h3339] = 8'h00;
mem[16'h333A] = 8'h00;
mem[16'h333B] = 8'h00;
mem[16'h333C] = 8'h00;
mem[16'h333D] = 8'h00;
mem[16'h333E] = 8'h00;
mem[16'h333F] = 8'h00;
mem[16'h3340] = 8'h00;
mem[16'h3341] = 8'h00;
mem[16'h3342] = 8'h00;
mem[16'h3343] = 8'h00;
mem[16'h3344] = 8'h00;
mem[16'h3345] = 8'h00;
mem[16'h3346] = 8'h00;
mem[16'h3347] = 8'h00;
mem[16'h3348] = 8'h00;
mem[16'h3349] = 8'h00;
mem[16'h334A] = 8'h00;
mem[16'h334B] = 8'h00;
mem[16'h334C] = 8'h00;
mem[16'h334D] = 8'h00;
mem[16'h334E] = 8'h00;
mem[16'h334F] = 8'h2A;
mem[16'h3350] = 8'h2A;
mem[16'h3351] = 8'h54;
mem[16'h3352] = 8'h0A;
mem[16'h3353] = 8'h55;
mem[16'h3354] = 8'h08;
mem[16'h3355] = 8'h55;
mem[16'h3356] = 8'h02;
mem[16'h3357] = 8'h41;
mem[16'h3358] = 8'h2A;
mem[16'h3359] = 8'h54;
mem[16'h335A] = 8'h0A;
mem[16'h335B] = 8'h55;
mem[16'h335C] = 8'h08;
mem[16'h335D] = 8'h55;
mem[16'h335E] = 8'h02;
mem[16'h335F] = 8'h41;
mem[16'h3360] = 8'h2A;
mem[16'h3361] = 8'h54;
mem[16'h3362] = 8'h60;
mem[16'h3363] = 8'h03;
mem[16'h3364] = 8'h08;
mem[16'h3365] = 8'h55;
mem[16'h3366] = 8'h02;
mem[16'h3367] = 8'h41;
mem[16'h3368] = 8'h2A;
mem[16'h3369] = 8'h54;
mem[16'h336A] = 8'h0A;
mem[16'h336B] = 8'h55;
mem[16'h336C] = 8'h08;
mem[16'h336D] = 8'h55;
mem[16'h336E] = 8'h02;
mem[16'h336F] = 8'h41;
mem[16'h3370] = 8'h2A;
mem[16'h3371] = 8'h54;
mem[16'h3372] = 8'h0A;
mem[16'h3373] = 8'h55;
mem[16'h3374] = 8'h08;
mem[16'h3375] = 8'h00;
mem[16'h3376] = 8'h00;
mem[16'h3377] = 8'h2A;
mem[16'h3378] = 8'h00;
mem[16'h3379] = 8'h00;
mem[16'h337A] = 8'h00;
mem[16'h337B] = 8'h00;
mem[16'h337C] = 8'h00;
mem[16'h337D] = 8'h00;
mem[16'h337E] = 8'h00;
mem[16'h337F] = 8'h00;
mem[16'h3380] = 8'hD5;
mem[16'h3381] = 8'hAA;
mem[16'h3382] = 8'hD5;
mem[16'h3383] = 8'hAA;
mem[16'h3384] = 8'hD5;
mem[16'h3385] = 8'hAA;
mem[16'h3386] = 8'hD5;
mem[16'h3387] = 8'hAA;
mem[16'h3388] = 8'hD5;
mem[16'h3389] = 8'hAA;
mem[16'h338A] = 8'hD5;
mem[16'h338B] = 8'hAA;
mem[16'h338C] = 8'hD5;
mem[16'h338D] = 8'hAA;
mem[16'h338E] = 8'hD5;
mem[16'h338F] = 8'hAA;
mem[16'h3390] = 8'hD5;
mem[16'h3391] = 8'hAA;
mem[16'h3392] = 8'hD5;
mem[16'h3393] = 8'hAA;
mem[16'h3394] = 8'hD5;
mem[16'h3395] = 8'hAA;
mem[16'h3396] = 8'hD5;
mem[16'h3397] = 8'hAA;
mem[16'h3398] = 8'hD5;
mem[16'h3399] = 8'hAA;
mem[16'h339A] = 8'hD5;
mem[16'h339B] = 8'hAA;
mem[16'h339C] = 8'hD5;
mem[16'h339D] = 8'hAA;
mem[16'h339E] = 8'hD5;
mem[16'h339F] = 8'hAA;
mem[16'h33A0] = 8'hD5;
mem[16'h33A1] = 8'hAA;
mem[16'h33A2] = 8'hD5;
mem[16'h33A3] = 8'hAA;
mem[16'h33A4] = 8'h85;
mem[16'h33A5] = 8'h00;
mem[16'h33A6] = 8'h00;
mem[16'h33A7] = 8'h00;
mem[16'h33A8] = 8'h00;
mem[16'h33A9] = 8'hA0;
mem[16'h33AA] = 8'h94;
mem[16'h33AB] = 8'h81;
mem[16'h33AC] = 8'h00;
mem[16'h33AD] = 8'h00;
mem[16'h33AE] = 8'h00;
mem[16'h33AF] = 8'h00;
mem[16'h33B0] = 8'h00;
mem[16'h33B1] = 8'h00;
mem[16'h33B2] = 8'h00;
mem[16'h33B3] = 8'h00;
mem[16'h33B4] = 8'h00;
mem[16'h33B5] = 8'h00;
mem[16'h33B6] = 8'h00;
mem[16'h33B7] = 8'h00;
mem[16'h33B8] = 8'h00;
mem[16'h33B9] = 8'h00;
mem[16'h33BA] = 8'h00;
mem[16'h33BB] = 8'h00;
mem[16'h33BC] = 8'h00;
mem[16'h33BD] = 8'h00;
mem[16'h33BE] = 8'h00;
mem[16'h33BF] = 8'h00;
mem[16'h33C0] = 8'h00;
mem[16'h33C1] = 8'h00;
mem[16'h33C2] = 8'h00;
mem[16'h33C3] = 8'h00;
mem[16'h33C4] = 8'h00;
mem[16'h33C5] = 8'h00;
mem[16'h33C6] = 8'h00;
mem[16'h33C7] = 8'h00;
mem[16'h33C8] = 8'h00;
mem[16'h33C9] = 8'h00;
mem[16'h33CA] = 8'h00;
mem[16'h33CB] = 8'h00;
mem[16'h33CC] = 8'h00;
mem[16'h33CD] = 8'h00;
mem[16'h33CE] = 8'h00;
mem[16'h33CF] = 8'h2A;
mem[16'h33D0] = 8'h22;
mem[16'h33D1] = 8'h15;
mem[16'h33D2] = 8'h22;
mem[16'h33D3] = 8'h55;
mem[16'h33D4] = 8'h20;
mem[16'h33D5] = 8'h50;
mem[16'h33D6] = 8'h0A;
mem[16'h33D7] = 8'h55;
mem[16'h33D8] = 8'h22;
mem[16'h33D9] = 8'h15;
mem[16'h33DA] = 8'h22;
mem[16'h33DB] = 8'h55;
mem[16'h33DC] = 8'h20;
mem[16'h33DD] = 8'h50;
mem[16'h33DE] = 8'h0A;
mem[16'h33DF] = 8'h55;
mem[16'h33E0] = 8'h22;
mem[16'h33E1] = 8'h15;
mem[16'h33E2] = 8'h22;
mem[16'h33E3] = 8'h55;
mem[16'h33E4] = 8'h20;
mem[16'h33E5] = 8'h50;
mem[16'h33E6] = 8'h0A;
mem[16'h33E7] = 8'h55;
mem[16'h33E8] = 8'h22;
mem[16'h33E9] = 8'h15;
mem[16'h33EA] = 8'h22;
mem[16'h33EB] = 8'h55;
mem[16'h33EC] = 8'h20;
mem[16'h33ED] = 8'h50;
mem[16'h33EE] = 8'h0A;
mem[16'h33EF] = 8'h55;
mem[16'h33F0] = 8'h22;
mem[16'h33F1] = 8'h15;
mem[16'h33F2] = 8'h22;
mem[16'h33F3] = 8'h55;
mem[16'h33F4] = 8'h00;
mem[16'h33F5] = 8'h62;
mem[16'h33F6] = 8'h00;
mem[16'h33F7] = 8'h2A;
mem[16'h33F8] = 8'h00;
mem[16'h33F9] = 8'h00;
mem[16'h33FA] = 8'h00;
mem[16'h33FB] = 8'h00;
mem[16'h33FC] = 8'h00;
mem[16'h33FD] = 8'h00;
mem[16'h33FE] = 8'h00;
mem[16'h33FF] = 8'h00;
mem[16'h3400] = 8'h00;
mem[16'h3401] = 8'h42;
mem[16'h3402] = 8'h10;
mem[16'h3403] = 8'h00;
mem[16'h3404] = 8'h42;
mem[16'h3405] = 8'h02;
mem[16'h3406] = 8'h44;
mem[16'h3407] = 8'h02;
mem[16'h3408] = 8'h02;
mem[16'h3409] = 8'h00;
mem[16'h340A] = 8'h42;
mem[16'h340B] = 8'h42;
mem[16'h340C] = 8'h42;
mem[16'h340D] = 8'h42;
mem[16'h340E] = 8'h42;
mem[16'h340F] = 8'h42;
mem[16'h3410] = 8'h00;
mem[16'h3411] = 8'h00;
mem[16'h3412] = 8'h00;
mem[16'h3413] = 8'h00;
mem[16'h3414] = 8'h10;
mem[16'h3415] = 8'h44;
mem[16'h3416] = 8'h62;
mem[16'h3417] = 8'h02;
mem[16'h3418] = 8'h00;
mem[16'h3419] = 8'h42;
mem[16'h341A] = 8'h02;
mem[16'h341B] = 8'h44;
mem[16'h341C] = 8'h02;
mem[16'h341D] = 8'h02;
mem[16'h341E] = 8'h00;
mem[16'h341F] = 8'h42;
mem[16'h3420] = 8'h42;
mem[16'h3421] = 8'h42;
mem[16'h3422] = 8'h42;
mem[16'h3423] = 8'h42;
mem[16'h3424] = 8'h42;
mem[16'h3425] = 8'h00;
mem[16'h3426] = 8'h60;
mem[16'h3427] = 8'h03;
mem[16'h3428] = 8'hD5;
mem[16'h3429] = 8'hAA;
mem[16'h342A] = 8'hD5;
mem[16'h342B] = 8'hAA;
mem[16'h342C] = 8'hB5;
mem[16'h342D] = 8'hD5;
mem[16'h342E] = 8'hAA;
mem[16'h342F] = 8'hD5;
mem[16'h3430] = 8'hAA;
mem[16'h3431] = 8'hD5;
mem[16'h3432] = 8'hAA;
mem[16'h3433] = 8'hD5;
mem[16'h3434] = 8'hD6;
mem[16'h3435] = 8'hAA;
mem[16'h3436] = 8'hD5;
mem[16'h3437] = 8'hAA;
mem[16'h3438] = 8'hD5;
mem[16'h3439] = 8'hD5;
mem[16'h343A] = 8'hAA;
mem[16'h343B] = 8'hD5;
mem[16'h343C] = 8'hAA;
mem[16'h343D] = 8'hD5;
mem[16'h343E] = 8'hAA;
mem[16'h343F] = 8'hD5;
mem[16'h3440] = 8'hDA;
mem[16'h3441] = 8'hAA;
mem[16'h3442] = 8'hD5;
mem[16'h3443] = 8'hAA;
mem[16'h3444] = 8'hAB;
mem[16'h3445] = 8'hD5;
mem[16'h3446] = 8'hAA;
mem[16'h3447] = 8'hD5;
mem[16'h3448] = 8'hAA;
mem[16'h3449] = 8'hD5;
mem[16'h344A] = 8'hAA;
mem[16'h344B] = 8'hB5;
mem[16'h344C] = 8'h85;
mem[16'h344D] = 8'h00;
mem[16'h344E] = 8'h00;
mem[16'h344F] = 8'h00;
mem[16'h3450] = 8'h00;
mem[16'h3451] = 8'h00;
mem[16'h3452] = 8'h00;
mem[16'h3453] = 8'h00;
mem[16'h3454] = 8'h00;
mem[16'h3455] = 8'h00;
mem[16'h3456] = 8'h00;
mem[16'h3457] = 8'h00;
mem[16'h3458] = 8'h00;
mem[16'h3459] = 8'h00;
mem[16'h345A] = 8'h00;
mem[16'h345B] = 8'h00;
mem[16'h345C] = 8'h00;
mem[16'h345D] = 8'h00;
mem[16'h345E] = 8'h00;
mem[16'h345F] = 8'h00;
mem[16'h3460] = 8'h00;
mem[16'h3461] = 8'h00;
mem[16'h3462] = 8'h00;
mem[16'h3463] = 8'h00;
mem[16'h3464] = 8'h00;
mem[16'h3465] = 8'h00;
mem[16'h3466] = 8'h00;
mem[16'h3467] = 8'h00;
mem[16'h3468] = 8'h00;
mem[16'h3469] = 8'h00;
mem[16'h346A] = 8'h00;
mem[16'h346B] = 8'h00;
mem[16'h346C] = 8'h00;
mem[16'h346D] = 8'h00;
mem[16'h346E] = 8'h00;
mem[16'h346F] = 8'h00;
mem[16'h3470] = 8'h00;
mem[16'h3471] = 8'h00;
mem[16'h3472] = 8'h00;
mem[16'h3473] = 8'h00;
mem[16'h3474] = 8'h00;
mem[16'h3475] = 8'h00;
mem[16'h3476] = 8'h00;
mem[16'h3477] = 8'h2A;
mem[16'h3478] = 8'h00;
mem[16'h3479] = 8'h00;
mem[16'h347A] = 8'h00;
mem[16'h347B] = 8'h00;
mem[16'h347C] = 8'h00;
mem[16'h347D] = 8'h00;
mem[16'h347E] = 8'h00;
mem[16'h347F] = 8'h00;
mem[16'h3480] = 8'h0A;
mem[16'h3481] = 8'h51;
mem[16'h3482] = 8'h2A;
mem[16'h3483] = 8'hAA;
mem[16'h3484] = 8'hD5;
mem[16'h3485] = 8'h45;
mem[16'h3486] = 8'h2A;
mem[16'h3487] = 8'h51;
mem[16'h3488] = 8'h0A;
mem[16'h3489] = 8'h51;
mem[16'h348A] = 8'hD5;
mem[16'h348B] = 8'hAA;
mem[16'h348C] = 8'h28;
mem[16'h348D] = 8'h45;
mem[16'h348E] = 8'h2A;
mem[16'h348F] = 8'h51;
mem[16'h3490] = 8'hD5;
mem[16'h3491] = 8'hAA;
mem[16'h3492] = 8'h2A;
mem[16'h3493] = 8'h10;
mem[16'h3494] = 8'h28;
mem[16'h3495] = 8'h45;
mem[16'h3496] = 8'h2A;
mem[16'h3497] = 8'hAA;
mem[16'h3498] = 8'hD5;
mem[16'h3499] = 8'h51;
mem[16'h349A] = 8'h2A;
mem[16'h349B] = 8'h10;
mem[16'h349C] = 8'h28;
mem[16'h349D] = 8'hAA;
mem[16'h349E] = 8'hD5;
mem[16'h349F] = 8'h51;
mem[16'h34A0] = 8'h0A;
mem[16'h34A1] = 8'h51;
mem[16'h34A2] = 8'h2A;
mem[16'h34A3] = 8'h10;
mem[16'h34A4] = 8'h08;
mem[16'h34A5] = 8'h00;
mem[16'h34A6] = 8'h0E;
mem[16'h34A7] = 8'h38;
mem[16'h34A8] = 8'hD5;
mem[16'h34A9] = 8'hAA;
mem[16'h34AA] = 8'hD5;
mem[16'h34AB] = 8'hAA;
mem[16'h34AC] = 8'hD5;
mem[16'h34AD] = 8'h8A;
mem[16'h34AE] = 8'hC5;
mem[16'h34AF] = 8'hAA;
mem[16'h34B0] = 8'hD1;
mem[16'h34B1] = 8'hA8;
mem[16'h34B2] = 8'h95;
mem[16'h34B3] = 8'h8A;
mem[16'h34B4] = 8'hD5;
mem[16'h34B5] = 8'hAA;
mem[16'h34B6] = 8'hD5;
mem[16'h34B7] = 8'hAA;
mem[16'h34B8] = 8'hD5;
mem[16'h34B9] = 8'hAA;
mem[16'h34BA] = 8'hD5;
mem[16'h34BB] = 8'hAA;
mem[16'h34BC] = 8'hC5;
mem[16'h34BD] = 8'hA2;
mem[16'h34BE] = 8'hD5;
mem[16'h34BF] = 8'hA8;
mem[16'h34C0] = 8'hD4;
mem[16'h34C1] = 8'h8A;
mem[16'h34C2] = 8'hC5;
mem[16'h34C3] = 8'hAA;
mem[16'h34C4] = 8'hD5;
mem[16'h34C5] = 8'hAA;
mem[16'h34C6] = 8'hD5;
mem[16'h34C7] = 8'hAA;
mem[16'h34C8] = 8'hD5;
mem[16'h34C9] = 8'hAA;
mem[16'h34CA] = 8'hD5;
mem[16'h34CB] = 8'hAA;
mem[16'h34CC] = 8'h85;
mem[16'h34CD] = 8'h00;
mem[16'h34CE] = 8'h00;
mem[16'h34CF] = 8'h2A;
mem[16'h34D0] = 8'h00;
mem[16'h34D1] = 8'h00;
mem[16'h34D2] = 8'h00;
mem[16'h34D3] = 8'h00;
mem[16'h34D4] = 8'h00;
mem[16'h34D5] = 8'h54;
mem[16'h34D6] = 8'h2A;
mem[16'h34D7] = 8'h03;
mem[16'h34D8] = 8'h00;
mem[16'h34D9] = 8'h00;
mem[16'h34DA] = 8'h00;
mem[16'h34DB] = 8'h00;
mem[16'h34DC] = 8'h00;
mem[16'h34DD] = 8'h00;
mem[16'h34DE] = 8'h00;
mem[16'h34DF] = 8'h00;
mem[16'h34E0] = 8'h00;
mem[16'h34E1] = 8'h54;
mem[16'h34E2] = 8'h2A;
mem[16'h34E3] = 8'h03;
mem[16'h34E4] = 8'h00;
mem[16'h34E5] = 8'h00;
mem[16'h34E6] = 8'h00;
mem[16'h34E7] = 8'h00;
mem[16'h34E8] = 8'h00;
mem[16'h34E9] = 8'h00;
mem[16'h34EA] = 8'h00;
mem[16'h34EB] = 8'h00;
mem[16'h34EC] = 8'h00;
mem[16'h34ED] = 8'h54;
mem[16'h34EE] = 8'h2A;
mem[16'h34EF] = 8'h03;
mem[16'h34F0] = 8'h00;
mem[16'h34F1] = 8'h00;
mem[16'h34F2] = 8'h00;
mem[16'h34F3] = 8'h00;
mem[16'h34F4] = 8'h00;
mem[16'h34F5] = 8'h00;
mem[16'h34F6] = 8'h00;
mem[16'h34F7] = 8'h2A;
mem[16'h34F8] = 8'h00;
mem[16'h34F9] = 8'h00;
mem[16'h34FA] = 8'h00;
mem[16'h34FB] = 8'h00;
mem[16'h34FC] = 8'h00;
mem[16'h34FD] = 8'h00;
mem[16'h34FE] = 8'h00;
mem[16'h34FF] = 8'h00;
mem[16'h3500] = 8'hD5;
mem[16'h3501] = 8'hAA;
mem[16'h3502] = 8'hD5;
mem[16'h3503] = 8'hAA;
mem[16'h3504] = 8'hD5;
mem[16'h3505] = 8'hAA;
mem[16'h3506] = 8'hD5;
mem[16'h3507] = 8'hAA;
mem[16'h3508] = 8'hD5;
mem[16'h3509] = 8'hAA;
mem[16'h350A] = 8'hD5;
mem[16'h350B] = 8'hAA;
mem[16'h350C] = 8'hD5;
mem[16'h350D] = 8'hAA;
mem[16'h350E] = 8'hD5;
mem[16'h350F] = 8'hAA;
mem[16'h3510] = 8'hD5;
mem[16'h3511] = 8'hAA;
mem[16'h3512] = 8'hD5;
mem[16'h3513] = 8'hAA;
mem[16'h3514] = 8'hD5;
mem[16'h3515] = 8'hAA;
mem[16'h3516] = 8'hD5;
mem[16'h3517] = 8'hAA;
mem[16'h3518] = 8'hD5;
mem[16'h3519] = 8'hAA;
mem[16'h351A] = 8'hD5;
mem[16'h351B] = 8'hAA;
mem[16'h351C] = 8'hD5;
mem[16'h351D] = 8'hAA;
mem[16'h351E] = 8'hD5;
mem[16'h351F] = 8'hAA;
mem[16'h3520] = 8'hD5;
mem[16'h3521] = 8'hAA;
mem[16'h3522] = 8'hD5;
mem[16'h3523] = 8'hAA;
mem[16'h3524] = 8'h85;
mem[16'h3525] = 8'h00;
mem[16'h3526] = 8'h60;
mem[16'h3527] = 8'h03;
mem[16'h3528] = 8'hD5;
mem[16'h3529] = 8'hAA;
mem[16'h352A] = 8'hD5;
mem[16'h352B] = 8'hAA;
mem[16'h352C] = 8'hD5;
mem[16'h352D] = 8'h8A;
mem[16'h352E] = 8'hC5;
mem[16'h352F] = 8'hAA;
mem[16'h3530] = 8'hD1;
mem[16'h3531] = 8'hA8;
mem[16'h3532] = 8'h95;
mem[16'h3533] = 8'h8A;
mem[16'h3534] = 8'hD5;
mem[16'h3535] = 8'hAA;
mem[16'h3536] = 8'hD5;
mem[16'h3537] = 8'hAA;
mem[16'h3538] = 8'hD5;
mem[16'h3539] = 8'hAA;
mem[16'h353A] = 8'hD5;
mem[16'h353B] = 8'hAA;
mem[16'h353C] = 8'hC5;
mem[16'h353D] = 8'hA2;
mem[16'h353E] = 8'hD5;
mem[16'h353F] = 8'hA8;
mem[16'h3540] = 8'hD4;
mem[16'h3541] = 8'h8A;
mem[16'h3542] = 8'hC5;
mem[16'h3543] = 8'hAA;
mem[16'h3544] = 8'hD5;
mem[16'h3545] = 8'hAA;
mem[16'h3546] = 8'hD5;
mem[16'h3547] = 8'hAA;
mem[16'h3548] = 8'hD5;
mem[16'h3549] = 8'hAA;
mem[16'h354A] = 8'hD5;
mem[16'h354B] = 8'hAA;
mem[16'h354C] = 8'h85;
mem[16'h354D] = 8'h00;
mem[16'h354E] = 8'h00;
mem[16'h354F] = 8'h2A;
mem[16'h3550] = 8'h00;
mem[16'h3551] = 8'hD8;
mem[16'h3552] = 8'h8D;
mem[16'h3553] = 8'h80;
mem[16'h3554] = 8'h00;
mem[16'h3555] = 8'h00;
mem[16'h3556] = 8'h00;
mem[16'h3557] = 8'h00;
mem[16'h3558] = 8'h00;
mem[16'h3559] = 8'h00;
mem[16'h355A] = 8'h00;
mem[16'h355B] = 8'hC0;
mem[16'h355C] = 8'hED;
mem[16'h355D] = 8'h80;
mem[16'h355E] = 8'h00;
mem[16'h355F] = 8'h00;
mem[16'h3560] = 8'h00;
mem[16'h3561] = 8'h00;
mem[16'h3562] = 8'h00;
mem[16'h3563] = 8'h00;
mem[16'h3564] = 8'h00;
mem[16'h3565] = 8'h00;
mem[16'h3566] = 8'hEC;
mem[16'h3567] = 8'h86;
mem[16'h3568] = 8'h80;
mem[16'h3569] = 8'h00;
mem[16'h356A] = 8'h00;
mem[16'h356B] = 8'h00;
mem[16'h356C] = 8'h00;
mem[16'h356D] = 8'h00;
mem[16'h356E] = 8'h00;
mem[16'h356F] = 8'h00;
mem[16'h3570] = 8'h00;
mem[16'h3571] = 8'h00;
mem[16'h3572] = 8'h00;
mem[16'h3573] = 8'h00;
mem[16'h3574] = 8'h00;
mem[16'h3575] = 8'h00;
mem[16'h3576] = 8'h00;
mem[16'h3577] = 8'h2A;
mem[16'h3578] = 8'h00;
mem[16'h3579] = 8'h00;
mem[16'h357A] = 8'h00;
mem[16'h357B] = 8'h00;
mem[16'h357C] = 8'h00;
mem[16'h357D] = 8'h00;
mem[16'h357E] = 8'h00;
mem[16'h357F] = 8'h00;
mem[16'h3580] = 8'hD5;
mem[16'h3581] = 8'hAA;
mem[16'h3582] = 8'hD5;
mem[16'h3583] = 8'hAA;
mem[16'h3584] = 8'hD5;
mem[16'h3585] = 8'hAA;
mem[16'h3586] = 8'hAB;
mem[16'h3587] = 8'hD5;
mem[16'h3588] = 8'hAA;
mem[16'h3589] = 8'hD5;
mem[16'h358A] = 8'hAA;
mem[16'h358B] = 8'hD5;
mem[16'h358C] = 8'hAA;
mem[16'h358D] = 8'hD5;
mem[16'h358E] = 8'hAA;
mem[16'h358F] = 8'hD5;
mem[16'h3590] = 8'hD5;
mem[16'h3591] = 8'hAA;
mem[16'h3592] = 8'hAD;
mem[16'h3593] = 8'hD5;
mem[16'h3594] = 8'hAA;
mem[16'h3595] = 8'hD5;
mem[16'h3596] = 8'hAA;
mem[16'h3597] = 8'hD5;
mem[16'h3598] = 8'hAA;
mem[16'h3599] = 8'hD5;
mem[16'h359A] = 8'hAA;
mem[16'h359B] = 8'hD5;
mem[16'h359C] = 8'hD6;
mem[16'h359D] = 8'hAA;
mem[16'h359E] = 8'hD5;
mem[16'h359F] = 8'hAA;
mem[16'h35A0] = 8'hD5;
mem[16'h35A1] = 8'hAA;
mem[16'h35A2] = 8'hD5;
mem[16'h35A3] = 8'hAA;
mem[16'h35A4] = 8'h85;
mem[16'h35A5] = 8'h00;
mem[16'h35A6] = 8'h00;
mem[16'h35A7] = 8'h00;
mem[16'h35A8] = 8'h02;
mem[16'h35A9] = 8'h55;
mem[16'h35AA] = 8'h28;
mem[16'h35AB] = 8'h15;
mem[16'h35AC] = 8'h2A;
mem[16'h35AD] = 8'h11;
mem[16'h35AE] = 8'h2A;
mem[16'h35AF] = 8'h05;
mem[16'h35B0] = 8'h02;
mem[16'h35B1] = 8'h55;
mem[16'h35B2] = 8'h28;
mem[16'h35B3] = 8'h15;
mem[16'h35B4] = 8'h2A;
mem[16'h35B5] = 8'h11;
mem[16'h35B6] = 8'h2A;
mem[16'h35B7] = 8'h05;
mem[16'h35B8] = 8'h02;
mem[16'h35B9] = 8'h55;
mem[16'h35BA] = 8'h28;
mem[16'h35BB] = 8'h15;
mem[16'h35BC] = 8'h2A;
mem[16'h35BD] = 8'h11;
mem[16'h35BE] = 8'h2A;
mem[16'h35BF] = 8'h05;
mem[16'h35C0] = 8'h02;
mem[16'h35C1] = 8'h55;
mem[16'h35C2] = 8'h28;
mem[16'h35C3] = 8'h15;
mem[16'h35C4] = 8'h2A;
mem[16'h35C5] = 8'h11;
mem[16'h35C6] = 8'h2A;
mem[16'h35C7] = 8'h05;
mem[16'h35C8] = 8'h02;
mem[16'h35C9] = 8'h55;
mem[16'h35CA] = 8'h28;
mem[16'h35CB] = 8'h15;
mem[16'h35CC] = 8'h0A;
mem[16'h35CD] = 8'h00;
mem[16'h35CE] = 8'h00;
mem[16'h35CF] = 8'h2A;
mem[16'h35D0] = 8'h00;
mem[16'h35D1] = 8'hD8;
mem[16'h35D2] = 8'h8D;
mem[16'h35D3] = 8'h80;
mem[16'h35D4] = 8'h00;
mem[16'h35D5] = 8'h00;
mem[16'h35D6] = 8'h00;
mem[16'h35D7] = 8'h00;
mem[16'h35D8] = 8'h00;
mem[16'h35D9] = 8'h00;
mem[16'h35DA] = 8'h00;
mem[16'h35DB] = 8'hC0;
mem[16'h35DC] = 8'hED;
mem[16'h35DD] = 8'h80;
mem[16'h35DE] = 8'h00;
mem[16'h35DF] = 8'h00;
mem[16'h35E0] = 8'h00;
mem[16'h35E1] = 8'h00;
mem[16'h35E2] = 8'h00;
mem[16'h35E3] = 8'h00;
mem[16'h35E4] = 8'h00;
mem[16'h35E5] = 8'h00;
mem[16'h35E6] = 8'hEC;
mem[16'h35E7] = 8'h86;
mem[16'h35E8] = 8'h80;
mem[16'h35E9] = 8'h00;
mem[16'h35EA] = 8'h00;
mem[16'h35EB] = 8'h00;
mem[16'h35EC] = 8'h00;
mem[16'h35ED] = 8'h00;
mem[16'h35EE] = 8'h00;
mem[16'h35EF] = 8'h00;
mem[16'h35F0] = 8'h00;
mem[16'h35F1] = 8'h00;
mem[16'h35F2] = 8'h00;
mem[16'h35F3] = 8'h00;
mem[16'h35F4] = 8'h00;
mem[16'h35F5] = 8'h00;
mem[16'h35F6] = 8'h00;
mem[16'h35F7] = 8'h2A;
mem[16'h35F8] = 8'h00;
mem[16'h35F9] = 8'h00;
mem[16'h35FA] = 8'h00;
mem[16'h35FB] = 8'h00;
mem[16'h35FC] = 8'h00;
mem[16'h35FD] = 8'h00;
mem[16'h35FE] = 8'h00;
mem[16'h35FF] = 8'h00;
mem[16'h3600] = 8'hD5;
mem[16'h3601] = 8'hA8;
mem[16'h3602] = 8'hD5;
mem[16'h3603] = 8'h8A;
mem[16'h3604] = 8'hD5;
mem[16'h3605] = 8'hAA;
mem[16'h3606] = 8'hD5;
mem[16'h3607] = 8'hAA;
mem[16'h3608] = 8'hD5;
mem[16'h3609] = 8'hA2;
mem[16'h360A] = 8'hD5;
mem[16'h360B] = 8'hAA;
mem[16'h360C] = 8'hD4;
mem[16'h360D] = 8'hAA;
mem[16'h360E] = 8'hD5;
mem[16'h360F] = 8'hAA;
mem[16'h3610] = 8'hD5;
mem[16'h3611] = 8'h8A;
mem[16'h3612] = 8'hD5;
mem[16'h3613] = 8'hAA;
mem[16'h3614] = 8'hD1;
mem[16'h3615] = 8'hAA;
mem[16'h3616] = 8'hD5;
mem[16'h3617] = 8'hAA;
mem[16'h3618] = 8'hD5;
mem[16'h3619] = 8'hAA;
mem[16'h361A] = 8'hD4;
mem[16'h361B] = 8'hAA;
mem[16'h361C] = 8'hC5;
mem[16'h361D] = 8'hAA;
mem[16'h361E] = 8'hD5;
mem[16'h361F] = 8'hAA;
mem[16'h3620] = 8'hD5;
mem[16'h3621] = 8'hAA;
mem[16'h3622] = 8'hD5;
mem[16'h3623] = 8'hAA;
mem[16'h3624] = 8'h85;
mem[16'h3625] = 8'h00;
mem[16'h3626] = 8'h74;
mem[16'h3627] = 8'h17;
mem[16'h3628] = 8'h02;
mem[16'h3629] = 8'h55;
mem[16'h362A] = 8'h28;
mem[16'h362B] = 8'h15;
mem[16'h362C] = 8'h2A;
mem[16'h362D] = 8'h11;
mem[16'h362E] = 8'h2A;
mem[16'h362F] = 8'h05;
mem[16'h3630] = 8'h02;
mem[16'h3631] = 8'h55;
mem[16'h3632] = 8'h28;
mem[16'h3633] = 8'h15;
mem[16'h3634] = 8'h2A;
mem[16'h3635] = 8'h11;
mem[16'h3636] = 8'h2A;
mem[16'h3637] = 8'h05;
mem[16'h3638] = 8'h02;
mem[16'h3639] = 8'h55;
mem[16'h363A] = 8'h28;
mem[16'h363B] = 8'h15;
mem[16'h363C] = 8'h2A;
mem[16'h363D] = 8'h11;
mem[16'h363E] = 8'h2A;
mem[16'h363F] = 8'h05;
mem[16'h3640] = 8'h02;
mem[16'h3641] = 8'h55;
mem[16'h3642] = 8'h28;
mem[16'h3643] = 8'h15;
mem[16'h3644] = 8'h2A;
mem[16'h3645] = 8'h11;
mem[16'h3646] = 8'h2A;
mem[16'h3647] = 8'h05;
mem[16'h3648] = 8'h02;
mem[16'h3649] = 8'h55;
mem[16'h364A] = 8'h28;
mem[16'h364B] = 8'h15;
mem[16'h364C] = 8'h0A;
mem[16'h364D] = 8'h00;
mem[16'h364E] = 8'h00;
mem[16'h364F] = 8'h2A;
mem[16'h3650] = 8'h00;
mem[16'h3651] = 8'h00;
mem[16'h3652] = 8'h00;
mem[16'h3653] = 8'h00;
mem[16'h3654] = 8'h56;
mem[16'h3655] = 8'h2A;
mem[16'h3656] = 8'h03;
mem[16'h3657] = 8'h00;
mem[16'h3658] = 8'h00;
mem[16'h3659] = 8'h00;
mem[16'h365A] = 8'h00;
mem[16'h365B] = 8'h00;
mem[16'h365C] = 8'h00;
mem[16'h365D] = 8'h00;
mem[16'h365E] = 8'h00;
mem[16'h365F] = 8'h00;
mem[16'h3660] = 8'h00;
mem[16'h3661] = 8'h00;
mem[16'h3662] = 8'h56;
mem[16'h3663] = 8'h2A;
mem[16'h3664] = 8'h03;
mem[16'h3665] = 8'h00;
mem[16'h3666] = 8'h00;
mem[16'h3667] = 8'h00;
mem[16'h3668] = 8'h00;
mem[16'h3669] = 8'h00;
mem[16'h366A] = 8'h00;
mem[16'h366B] = 8'h00;
mem[16'h366C] = 8'h00;
mem[16'h366D] = 8'h00;
mem[16'h366E] = 8'h00;
mem[16'h366F] = 8'h00;
mem[16'h3670] = 8'h56;
mem[16'h3671] = 8'h2A;
mem[16'h3672] = 8'h03;
mem[16'h3673] = 8'h00;
mem[16'h3674] = 8'h00;
mem[16'h3675] = 8'h00;
mem[16'h3676] = 8'h00;
mem[16'h3677] = 8'h2A;
mem[16'h3678] = 8'h00;
mem[16'h3679] = 8'h00;
mem[16'h367A] = 8'h00;
mem[16'h367B] = 8'h00;
mem[16'h367C] = 8'h00;
mem[16'h367D] = 8'h00;
mem[16'h367E] = 8'h00;
mem[16'h367F] = 8'h00;
mem[16'h3680] = 8'hD5;
mem[16'h3681] = 8'h94;
mem[16'h3682] = 8'hD4;
mem[16'h3683] = 8'hCA;
mem[16'h3684] = 8'hC2;
mem[16'h3685] = 8'hAA;
mem[16'h3686] = 8'hD5;
mem[16'h3687] = 8'hAA;
mem[16'h3688] = 8'hD5;
mem[16'h3689] = 8'hD2;
mem[16'h368A] = 8'hD0;
mem[16'h368B] = 8'hAA;
mem[16'h368C] = 8'h8A;
mem[16'h368D] = 8'hAA;
mem[16'h368E] = 8'hD5;
mem[16'h368F] = 8'hAA;
mem[16'h3690] = 8'hD5;
mem[16'h3691] = 8'hCA;
mem[16'h3692] = 8'hC2;
mem[16'h3693] = 8'hAA;
mem[16'h3694] = 8'hA9;
mem[16'h3695] = 8'hA8;
mem[16'h3696] = 8'hD5;
mem[16'h3697] = 8'hAA;
mem[16'h3698] = 8'hD5;
mem[16'h3699] = 8'hAA;
mem[16'h369A] = 8'h8A;
mem[16'h369B] = 8'hAA;
mem[16'h369C] = 8'hA5;
mem[16'h369D] = 8'hA1;
mem[16'h369E] = 8'hD5;
mem[16'h369F] = 8'hAA;
mem[16'h36A0] = 8'hD5;
mem[16'h36A1] = 8'hAA;
mem[16'h36A2] = 8'hD5;
mem[16'h36A3] = 8'hAA;
mem[16'h36A4] = 8'h85;
mem[16'h36A5] = 8'h00;
mem[16'h36A6] = 8'h40;
mem[16'h36A7] = 8'h01;
mem[16'h36A8] = 8'h00;
mem[16'h36A9] = 8'h00;
mem[16'h36AA] = 8'h1E;
mem[16'h36AB] = 8'h55;
mem[16'h36AC] = 8'h0A;
mem[16'h36AD] = 8'h00;
mem[16'h36AE] = 8'h00;
mem[16'h36AF] = 8'h00;
mem[16'h36B0] = 8'h00;
mem[16'h36B1] = 8'h00;
mem[16'h36B2] = 8'h00;
mem[16'h36B3] = 8'h00;
mem[16'h36B4] = 8'h00;
mem[16'h36B5] = 8'h00;
mem[16'h36B6] = 8'h00;
mem[16'h36B7] = 8'h00;
mem[16'h36B8] = 8'h1E;
mem[16'h36B9] = 8'h55;
mem[16'h36BA] = 8'h0A;
mem[16'h36BB] = 8'h00;
mem[16'h36BC] = 8'h00;
mem[16'h36BD] = 8'h00;
mem[16'h36BE] = 8'h00;
mem[16'h36BF] = 8'h00;
mem[16'h36C0] = 8'h00;
mem[16'h36C1] = 8'h00;
mem[16'h36C2] = 8'h00;
mem[16'h36C3] = 8'h00;
mem[16'h36C4] = 8'h00;
mem[16'h36C5] = 8'h00;
mem[16'h36C6] = 8'h00;
mem[16'h36C7] = 8'h00;
mem[16'h36C8] = 8'h00;
mem[16'h36C9] = 8'h00;
mem[16'h36CA] = 8'h00;
mem[16'h36CB] = 8'h00;
mem[16'h36CC] = 8'h00;
mem[16'h36CD] = 8'h00;
mem[16'h36CE] = 8'h00;
mem[16'h36CF] = 8'h2A;
mem[16'h36D0] = 8'h00;
mem[16'h36D1] = 8'h00;
mem[16'h36D2] = 8'h00;
mem[16'h36D3] = 8'h00;
mem[16'h36D4] = 8'h00;
mem[16'h36D5] = 8'h00;
mem[16'h36D6] = 8'h00;
mem[16'h36D7] = 8'h00;
mem[16'h36D8] = 8'h00;
mem[16'h36D9] = 8'h00;
mem[16'h36DA] = 8'h00;
mem[16'h36DB] = 8'h00;
mem[16'h36DC] = 8'h00;
mem[16'h36DD] = 8'h00;
mem[16'h36DE] = 8'h00;
mem[16'h36DF] = 8'h00;
mem[16'h36E0] = 8'h00;
mem[16'h36E1] = 8'h00;
mem[16'h36E2] = 8'h00;
mem[16'h36E3] = 8'h00;
mem[16'h36E4] = 8'h00;
mem[16'h36E5] = 8'h00;
mem[16'h36E6] = 8'h00;
mem[16'h36E7] = 8'h00;
mem[16'h36E8] = 8'h00;
mem[16'h36E9] = 8'h00;
mem[16'h36EA] = 8'h00;
mem[16'h36EB] = 8'h00;
mem[16'h36EC] = 8'h00;
mem[16'h36ED] = 8'h00;
mem[16'h36EE] = 8'h00;
mem[16'h36EF] = 8'h00;
mem[16'h36F0] = 8'h00;
mem[16'h36F1] = 8'h00;
mem[16'h36F2] = 8'h00;
mem[16'h36F3] = 8'h00;
mem[16'h36F4] = 8'h00;
mem[16'h36F5] = 8'h00;
mem[16'h36F6] = 8'h00;
mem[16'h36F7] = 8'h2A;
mem[16'h36F8] = 8'h00;
mem[16'h36F9] = 8'h00;
mem[16'h36FA] = 8'h00;
mem[16'h36FB] = 8'h00;
mem[16'h36FC] = 8'h00;
mem[16'h36FD] = 8'h00;
mem[16'h36FE] = 8'h00;
mem[16'h36FF] = 8'h00;
mem[16'h3700] = 8'hAB;
mem[16'h3701] = 8'hAD;
mem[16'h3702] = 8'hD5;
mem[16'h3703] = 8'hAA;
mem[16'h3704] = 8'hD5;
mem[16'h3705] = 8'hAA;
mem[16'h3706] = 8'hD5;
mem[16'h3707] = 8'hAA;
mem[16'h3708] = 8'hD5;
mem[16'h3709] = 8'hAA;
mem[16'h370A] = 8'hD5;
mem[16'h370B] = 8'hD5;
mem[16'h370C] = 8'hAA;
mem[16'h370D] = 8'hD5;
mem[16'h370E] = 8'hAA;
mem[16'h370F] = 8'hD5;
mem[16'h3710] = 8'hAA;
mem[16'h3711] = 8'hD5;
mem[16'h3712] = 8'hAA;
mem[16'h3713] = 8'hD5;
mem[16'h3714] = 8'hAA;
mem[16'h3715] = 8'hD5;
mem[16'h3716] = 8'hAA;
mem[16'h3717] = 8'hD5;
mem[16'h3718] = 8'hAA;
mem[16'h3719] = 8'hD5;
mem[16'h371A] = 8'hD5;
mem[16'h371B] = 8'hAA;
mem[16'h371C] = 8'hD5;
mem[16'h371D] = 8'hAA;
mem[16'h371E] = 8'hD5;
mem[16'h371F] = 8'hAA;
mem[16'h3720] = 8'hD5;
mem[16'h3721] = 8'hAA;
mem[16'h3722] = 8'hD5;
mem[16'h3723] = 8'hAA;
mem[16'h3724] = 8'h85;
mem[16'h3725] = 8'h00;
mem[16'h3726] = 8'h7C;
mem[16'h3727] = 8'h1F;
mem[16'h3728] = 8'h00;
mem[16'h3729] = 8'h00;
mem[16'h372A] = 8'h00;
mem[16'h372B] = 8'h00;
mem[16'h372C] = 8'h00;
mem[16'h372D] = 8'h00;
mem[16'h372E] = 8'h00;
mem[16'h372F] = 8'h00;
mem[16'h3730] = 8'h00;
mem[16'h3731] = 8'h00;
mem[16'h3732] = 8'h00;
mem[16'h3733] = 8'h00;
mem[16'h3734] = 8'h00;
mem[16'h3735] = 8'h00;
mem[16'h3736] = 8'h00;
mem[16'h3737] = 8'h00;
mem[16'h3738] = 8'h00;
mem[16'h3739] = 8'h00;
mem[16'h373A] = 8'h00;
mem[16'h373B] = 8'h00;
mem[16'h373C] = 8'h00;
mem[16'h373D] = 8'h00;
mem[16'h373E] = 8'h00;
mem[16'h373F] = 8'h00;
mem[16'h3740] = 8'h00;
mem[16'h3741] = 8'h00;
mem[16'h3742] = 8'h00;
mem[16'h3743] = 8'h00;
mem[16'h3744] = 8'h00;
mem[16'h3745] = 8'h00;
mem[16'h3746] = 8'h00;
mem[16'h3747] = 8'h00;
mem[16'h3748] = 8'h00;
mem[16'h3749] = 8'h00;
mem[16'h374A] = 8'h00;
mem[16'h374B] = 8'h00;
mem[16'h374C] = 8'h00;
mem[16'h374D] = 8'h00;
mem[16'h374E] = 8'h00;
mem[16'h374F] = 8'h2A;
mem[16'h3750] = 8'h28;
mem[16'h3751] = 8'h15;
mem[16'h3752] = 8'h08;
mem[16'h3753] = 8'h54;
mem[16'h3754] = 8'h22;
mem[16'h3755] = 8'h55;
mem[16'h3756] = 8'h28;
mem[16'h3757] = 8'h45;
mem[16'h3758] = 8'h28;
mem[16'h3759] = 8'h15;
mem[16'h375A] = 8'h08;
mem[16'h375B] = 8'h54;
mem[16'h375C] = 8'h22;
mem[16'h375D] = 8'h55;
mem[16'h375E] = 8'h28;
mem[16'h375F] = 8'h45;
mem[16'h3760] = 8'h28;
mem[16'h3761] = 8'h15;
mem[16'h3762] = 8'h70;
mem[16'h3763] = 8'h07;
mem[16'h3764] = 8'h22;
mem[16'h3765] = 8'h55;
mem[16'h3766] = 8'h28;
mem[16'h3767] = 8'h45;
mem[16'h3768] = 8'h28;
mem[16'h3769] = 8'h15;
mem[16'h376A] = 8'h08;
mem[16'h376B] = 8'h54;
mem[16'h376C] = 8'h22;
mem[16'h376D] = 8'h55;
mem[16'h376E] = 8'h28;
mem[16'h376F] = 8'h45;
mem[16'h3770] = 8'h28;
mem[16'h3771] = 8'h15;
mem[16'h3772] = 8'h08;
mem[16'h3773] = 8'h54;
mem[16'h3774] = 8'h02;
mem[16'h3775] = 8'h00;
mem[16'h3776] = 8'h00;
mem[16'h3777] = 8'h2A;
mem[16'h3778] = 8'h00;
mem[16'h3779] = 8'h00;
mem[16'h377A] = 8'h00;
mem[16'h377B] = 8'h00;
mem[16'h377C] = 8'h00;
mem[16'h377D] = 8'h00;
mem[16'h377E] = 8'h00;
mem[16'h377F] = 8'h00;
mem[16'h3780] = 8'hD5;
mem[16'h3781] = 8'hAA;
mem[16'h3782] = 8'hD5;
mem[16'h3783] = 8'hAA;
mem[16'h3784] = 8'hD5;
mem[16'h3785] = 8'hAA;
mem[16'h3786] = 8'hD5;
mem[16'h3787] = 8'hAA;
mem[16'h3788] = 8'hD5;
mem[16'h3789] = 8'hAA;
mem[16'h378A] = 8'hD5;
mem[16'h378B] = 8'hAA;
mem[16'h378C] = 8'hD5;
mem[16'h378D] = 8'hAA;
mem[16'h378E] = 8'hD5;
mem[16'h378F] = 8'hAA;
mem[16'h3790] = 8'hD5;
mem[16'h3791] = 8'hAA;
mem[16'h3792] = 8'hD5;
mem[16'h3793] = 8'hAA;
mem[16'h3794] = 8'hD5;
mem[16'h3795] = 8'hAA;
mem[16'h3796] = 8'hD5;
mem[16'h3797] = 8'hAA;
mem[16'h3798] = 8'hD5;
mem[16'h3799] = 8'hAA;
mem[16'h379A] = 8'hD5;
mem[16'h379B] = 8'hAA;
mem[16'h379C] = 8'hD5;
mem[16'h379D] = 8'hAA;
mem[16'h379E] = 8'hD5;
mem[16'h379F] = 8'hAA;
mem[16'h37A0] = 8'hD5;
mem[16'h37A1] = 8'hAA;
mem[16'h37A2] = 8'hD5;
mem[16'h37A3] = 8'hAA;
mem[16'h37A4] = 8'h85;
mem[16'h37A5] = 8'h00;
mem[16'h37A6] = 8'h00;
mem[16'h37A7] = 8'h00;
mem[16'h37A8] = 8'h00;
mem[16'h37A9] = 8'hA0;
mem[16'h37AA] = 8'hD5;
mem[16'h37AB] = 8'h82;
mem[16'h37AC] = 8'h00;
mem[16'h37AD] = 8'h00;
mem[16'h37AE] = 8'h00;
mem[16'h37AF] = 8'h00;
mem[16'h37B0] = 8'h00;
mem[16'h37B1] = 8'h00;
mem[16'h37B2] = 8'h00;
mem[16'h37B3] = 8'h00;
mem[16'h37B4] = 8'h00;
mem[16'h37B5] = 8'h00;
mem[16'h37B6] = 8'h00;
mem[16'h37B7] = 8'h00;
mem[16'h37B8] = 8'h00;
mem[16'h37B9] = 8'h00;
mem[16'h37BA] = 8'h00;
mem[16'h37BB] = 8'h00;
mem[16'h37BC] = 8'h00;
mem[16'h37BD] = 8'h00;
mem[16'h37BE] = 8'h00;
mem[16'h37BF] = 8'h00;
mem[16'h37C0] = 8'h00;
mem[16'h37C1] = 8'h00;
mem[16'h37C2] = 8'h00;
mem[16'h37C3] = 8'h00;
mem[16'h37C4] = 8'h00;
mem[16'h37C5] = 8'h00;
mem[16'h37C6] = 8'h00;
mem[16'h37C7] = 8'h00;
mem[16'h37C8] = 8'h00;
mem[16'h37C9] = 8'h00;
mem[16'h37CA] = 8'h00;
mem[16'h37CB] = 8'h00;
mem[16'h37CC] = 8'h00;
mem[16'h37CD] = 8'h00;
mem[16'h37CE] = 8'h00;
mem[16'h37CF] = 8'h2A;
mem[16'h37D0] = 8'h02;
mem[16'h37D1] = 8'h55;
mem[16'h37D2] = 8'h28;
mem[16'h37D3] = 8'h15;
mem[16'h37D4] = 8'h2A;
mem[16'h37D5] = 8'h11;
mem[16'h37D6] = 8'h2A;
mem[16'h37D7] = 8'h05;
mem[16'h37D8] = 8'h02;
mem[16'h37D9] = 8'h55;
mem[16'h37DA] = 8'h28;
mem[16'h37DB] = 8'h15;
mem[16'h37DC] = 8'h2A;
mem[16'h37DD] = 8'h11;
mem[16'h37DE] = 8'h2A;
mem[16'h37DF] = 8'h05;
mem[16'h37E0] = 8'h02;
mem[16'h37E1] = 8'h55;
mem[16'h37E2] = 8'h28;
mem[16'h37E3] = 8'h15;
mem[16'h37E4] = 8'h2A;
mem[16'h37E5] = 8'h11;
mem[16'h37E6] = 8'h2A;
mem[16'h37E7] = 8'h05;
mem[16'h37E8] = 8'h02;
mem[16'h37E9] = 8'h55;
mem[16'h37EA] = 8'h28;
mem[16'h37EB] = 8'h15;
mem[16'h37EC] = 8'h2A;
mem[16'h37ED] = 8'h11;
mem[16'h37EE] = 8'h2A;
mem[16'h37EF] = 8'h05;
mem[16'h37F0] = 8'h02;
mem[16'h37F1] = 8'h55;
mem[16'h37F2] = 8'h28;
mem[16'h37F3] = 8'h15;
mem[16'h37F4] = 8'h0A;
mem[16'h37F5] = 8'h42;
mem[16'h37F6] = 8'h00;
mem[16'h37F7] = 8'h2A;
mem[16'h37F8] = 8'h00;
mem[16'h37F9] = 8'h00;
mem[16'h37FA] = 8'h00;
mem[16'h37FB] = 8'h00;
mem[16'h37FC] = 8'h00;
mem[16'h37FD] = 8'h00;
mem[16'h37FE] = 8'h00;
mem[16'h37FF] = 8'h00;
mem[16'h3800] = 8'h00;
mem[16'h3801] = 8'h42;
mem[16'h3802] = 8'h38;
mem[16'h3803] = 8'h00;
mem[16'h3804] = 8'h3C;
mem[16'h3805] = 8'h3C;
mem[16'h3806] = 8'h38;
mem[16'h3807] = 8'h02;
mem[16'h3808] = 8'h3C;
mem[16'h3809] = 8'h00;
mem[16'h380A] = 8'h3C;
mem[16'h380B] = 8'h3C;
mem[16'h380C] = 8'h3C;
mem[16'h380D] = 8'h3C;
mem[16'h380E] = 8'h3C;
mem[16'h380F] = 8'h3C;
mem[16'h3810] = 8'h00;
mem[16'h3811] = 8'h00;
mem[16'h3812] = 8'h00;
mem[16'h3813] = 8'h00;
mem[16'h3814] = 8'h10;
mem[16'h3815] = 8'h38;
mem[16'h3816] = 8'h5C;
mem[16'h3817] = 8'h02;
mem[16'h3818] = 8'h00;
mem[16'h3819] = 8'h3C;
mem[16'h381A] = 8'h3C;
mem[16'h381B] = 8'h38;
mem[16'h381C] = 8'h02;
mem[16'h381D] = 8'h3C;
mem[16'h381E] = 8'h00;
mem[16'h381F] = 8'h3C;
mem[16'h3820] = 8'h3C;
mem[16'h3821] = 8'h3C;
mem[16'h3822] = 8'h3C;
mem[16'h3823] = 8'h3C;
mem[16'h3824] = 8'h3C;
mem[16'h3825] = 8'h00;
mem[16'h3826] = 8'h40;
mem[16'h3827] = 8'h01;
mem[16'h3828] = 8'hD5;
mem[16'h3829] = 8'hAA;
mem[16'h382A] = 8'hD5;
mem[16'h382B] = 8'hAA;
mem[16'h382C] = 8'hB5;
mem[16'h382D] = 8'hD5;
mem[16'h382E] = 8'hAA;
mem[16'h382F] = 8'hD5;
mem[16'h3830] = 8'hAA;
mem[16'h3831] = 8'hD5;
mem[16'h3832] = 8'hAA;
mem[16'h3833] = 8'hD5;
mem[16'h3834] = 8'hD6;
mem[16'h3835] = 8'hAA;
mem[16'h3836] = 8'hD5;
mem[16'h3837] = 8'hAA;
mem[16'h3838] = 8'hD5;
mem[16'h3839] = 8'hD5;
mem[16'h383A] = 8'hAA;
mem[16'h383B] = 8'hD5;
mem[16'h383C] = 8'hAA;
mem[16'h383D] = 8'hD5;
mem[16'h383E] = 8'hAA;
mem[16'h383F] = 8'hD5;
mem[16'h3840] = 8'hDA;
mem[16'h3841] = 8'hAA;
mem[16'h3842] = 8'hD5;
mem[16'h3843] = 8'hAA;
mem[16'h3844] = 8'hAB;
mem[16'h3845] = 8'hD5;
mem[16'h3846] = 8'hAA;
mem[16'h3847] = 8'hD5;
mem[16'h3848] = 8'hAA;
mem[16'h3849] = 8'hD5;
mem[16'h384A] = 8'hAA;
mem[16'h384B] = 8'hB5;
mem[16'h384C] = 8'h85;
mem[16'h384D] = 8'h00;
mem[16'h384E] = 8'h00;
mem[16'h384F] = 8'h2A;
mem[16'h3850] = 8'h00;
mem[16'h3851] = 8'h00;
mem[16'h3852] = 8'h00;
mem[16'h3853] = 8'h00;
mem[16'h3854] = 8'h00;
mem[16'h3855] = 8'h00;
mem[16'h3856] = 8'h00;
mem[16'h3857] = 8'h00;
mem[16'h3858] = 8'h00;
mem[16'h3859] = 8'h00;
mem[16'h385A] = 8'h00;
mem[16'h385B] = 8'h00;
mem[16'h385C] = 8'h00;
mem[16'h385D] = 8'h00;
mem[16'h385E] = 8'h00;
mem[16'h385F] = 8'h00;
mem[16'h3860] = 8'h00;
mem[16'h3861] = 8'h00;
mem[16'h3862] = 8'h00;
mem[16'h3863] = 8'h00;
mem[16'h3864] = 8'h00;
mem[16'h3865] = 8'h00;
mem[16'h3866] = 8'h00;
mem[16'h3867] = 8'h00;
mem[16'h3868] = 8'h00;
mem[16'h3869] = 8'h00;
mem[16'h386A] = 8'h00;
mem[16'h386B] = 8'h00;
mem[16'h386C] = 8'h00;
mem[16'h386D] = 8'h00;
mem[16'h386E] = 8'h00;
mem[16'h386F] = 8'h00;
mem[16'h3870] = 8'h00;
mem[16'h3871] = 8'h00;
mem[16'h3872] = 8'h00;
mem[16'h3873] = 8'h00;
mem[16'h3874] = 8'h00;
mem[16'h3875] = 8'h00;
mem[16'h3876] = 8'h00;
mem[16'h3877] = 8'h2A;
mem[16'h3878] = 8'h00;
mem[16'h3879] = 8'h00;
mem[16'h387A] = 8'h00;
mem[16'h387B] = 8'h00;
mem[16'h387C] = 8'h00;
mem[16'h387D] = 8'h00;
mem[16'h387E] = 8'h00;
mem[16'h387F] = 8'h00;
mem[16'h3880] = 8'h2A;
mem[16'h3881] = 8'h54;
mem[16'h3882] = 8'h0A;
mem[16'h3883] = 8'hAA;
mem[16'h3884] = 8'hD5;
mem[16'h3885] = 8'h55;
mem[16'h3886] = 8'h02;
mem[16'h3887] = 8'h41;
mem[16'h3888] = 8'h2A;
mem[16'h3889] = 8'h54;
mem[16'h388A] = 8'hD5;
mem[16'h388B] = 8'hAA;
mem[16'h388C] = 8'h08;
mem[16'h388D] = 8'h55;
mem[16'h388E] = 8'h02;
mem[16'h388F] = 8'h41;
mem[16'h3890] = 8'hD5;
mem[16'h3891] = 8'hAA;
mem[16'h3892] = 8'h0A;
mem[16'h3893] = 8'h55;
mem[16'h3894] = 8'h08;
mem[16'h3895] = 8'h55;
mem[16'h3896] = 8'h02;
mem[16'h3897] = 8'hAA;
mem[16'h3898] = 8'hD5;
mem[16'h3899] = 8'h54;
mem[16'h389A] = 8'h0A;
mem[16'h389B] = 8'h55;
mem[16'h389C] = 8'h08;
mem[16'h389D] = 8'hAA;
mem[16'h389E] = 8'hD5;
mem[16'h389F] = 8'h41;
mem[16'h38A0] = 8'h2A;
mem[16'h38A1] = 8'h54;
mem[16'h38A2] = 8'h0A;
mem[16'h38A3] = 8'h55;
mem[16'h38A4] = 8'h08;
mem[16'h38A5] = 8'h00;
mem[16'h38A6] = 8'h0E;
mem[16'h38A7] = 8'h38;
mem[16'h38A8] = 8'hD5;
mem[16'h38A9] = 8'hAA;
mem[16'h38AA] = 8'hD5;
mem[16'h38AB] = 8'hAA;
mem[16'h38AC] = 8'hD5;
mem[16'h38AD] = 8'hCA;
mem[16'h38AE] = 8'hC2;
mem[16'h38AF] = 8'hAA;
mem[16'h38B0] = 8'hA9;
mem[16'h38B1] = 8'hA8;
mem[16'h38B2] = 8'h95;
mem[16'h38B3] = 8'h85;
mem[16'h38B4] = 8'hD5;
mem[16'h38B5] = 8'hAA;
mem[16'h38B6] = 8'hD5;
mem[16'h38B7] = 8'hAA;
mem[16'h38B8] = 8'hD5;
mem[16'h38B9] = 8'hAA;
mem[16'h38BA] = 8'hD5;
mem[16'h38BB] = 8'hAA;
mem[16'h38BC] = 8'hA5;
mem[16'h38BD] = 8'hA1;
mem[16'h38BE] = 8'hD5;
mem[16'h38BF] = 8'h94;
mem[16'h38C0] = 8'hD4;
mem[16'h38C1] = 8'hCA;
mem[16'h38C2] = 8'hC2;
mem[16'h38C3] = 8'hAA;
mem[16'h38C4] = 8'hD5;
mem[16'h38C5] = 8'hAA;
mem[16'h38C6] = 8'hD5;
mem[16'h38C7] = 8'hAA;
mem[16'h38C8] = 8'hD5;
mem[16'h38C9] = 8'hAA;
mem[16'h38CA] = 8'hD5;
mem[16'h38CB] = 8'hAA;
mem[16'h38CC] = 8'h85;
mem[16'h38CD] = 8'h00;
mem[16'h38CE] = 8'h00;
mem[16'h38CF] = 8'h2A;
mem[16'h38D0] = 8'h00;
mem[16'h38D1] = 8'h00;
mem[16'h38D2] = 8'h00;
mem[16'h38D3] = 8'h00;
mem[16'h38D4] = 8'h00;
mem[16'h38D5] = 8'h78;
mem[16'h38D6] = 8'h30;
mem[16'h38D7] = 8'h01;
mem[16'h38D8] = 8'h00;
mem[16'h38D9] = 8'h00;
mem[16'h38DA] = 8'h00;
mem[16'h38DB] = 8'h00;
mem[16'h38DC] = 8'h00;
mem[16'h38DD] = 8'h00;
mem[16'h38DE] = 8'h00;
mem[16'h38DF] = 8'h00;
mem[16'h38E0] = 8'h00;
mem[16'h38E1] = 8'h78;
mem[16'h38E2] = 8'h30;
mem[16'h38E3] = 8'h01;
mem[16'h38E4] = 8'h00;
mem[16'h38E5] = 8'h00;
mem[16'h38E6] = 8'h00;
mem[16'h38E7] = 8'h00;
mem[16'h38E8] = 8'h00;
mem[16'h38E9] = 8'h00;
mem[16'h38EA] = 8'h00;
mem[16'h38EB] = 8'h00;
mem[16'h38EC] = 8'h00;
mem[16'h38ED] = 8'h78;
mem[16'h38EE] = 8'h30;
mem[16'h38EF] = 8'h01;
mem[16'h38F0] = 8'h00;
mem[16'h38F1] = 8'h00;
mem[16'h38F2] = 8'h00;
mem[16'h38F3] = 8'h00;
mem[16'h38F4] = 8'h00;
mem[16'h38F5] = 8'h00;
mem[16'h38F6] = 8'h00;
mem[16'h38F7] = 8'h2A;
mem[16'h38F8] = 8'h00;
mem[16'h38F9] = 8'h00;
mem[16'h38FA] = 8'h00;
mem[16'h38FB] = 8'h00;
mem[16'h38FC] = 8'h00;
mem[16'h38FD] = 8'h00;
mem[16'h38FE] = 8'h00;
mem[16'h38FF] = 8'h00;
mem[16'h3900] = 8'hD5;
mem[16'h3901] = 8'hAA;
mem[16'h3902] = 8'hD5;
mem[16'h3903] = 8'hAA;
mem[16'h3904] = 8'hD5;
mem[16'h3905] = 8'hAA;
mem[16'h3906] = 8'hD5;
mem[16'h3907] = 8'hAA;
mem[16'h3908] = 8'hD5;
mem[16'h3909] = 8'hAA;
mem[16'h390A] = 8'hD5;
mem[16'h390B] = 8'hAA;
mem[16'h390C] = 8'hD5;
mem[16'h390D] = 8'hAA;
mem[16'h390E] = 8'hD5;
mem[16'h390F] = 8'hAA;
mem[16'h3910] = 8'hD5;
mem[16'h3911] = 8'hAA;
mem[16'h3912] = 8'hD5;
mem[16'h3913] = 8'hAA;
mem[16'h3914] = 8'hD5;
mem[16'h3915] = 8'hAA;
mem[16'h3916] = 8'hD5;
mem[16'h3917] = 8'hAA;
mem[16'h3918] = 8'hD5;
mem[16'h3919] = 8'hAA;
mem[16'h391A] = 8'hD5;
mem[16'h391B] = 8'hAA;
mem[16'h391C] = 8'hD5;
mem[16'h391D] = 8'hAA;
mem[16'h391E] = 8'hD5;
mem[16'h391F] = 8'hAA;
mem[16'h3920] = 8'hD5;
mem[16'h3921] = 8'hAA;
mem[16'h3922] = 8'hD5;
mem[16'h3923] = 8'hAA;
mem[16'h3924] = 8'h85;
mem[16'h3925] = 8'h00;
mem[16'h3926] = 8'h70;
mem[16'h3927] = 8'h07;
mem[16'h3928] = 8'hD5;
mem[16'h3929] = 8'hAA;
mem[16'h392A] = 8'hD5;
mem[16'h392B] = 8'hAA;
mem[16'h392C] = 8'hD5;
mem[16'h392D] = 8'h8A;
mem[16'h392E] = 8'hD5;
mem[16'h392F] = 8'hAA;
mem[16'h3930] = 8'hD1;
mem[16'h3931] = 8'hAA;
mem[16'h3932] = 8'h95;
mem[16'h3933] = 8'hAA;
mem[16'h3934] = 8'hD5;
mem[16'h3935] = 8'hAA;
mem[16'h3936] = 8'hD5;
mem[16'h3937] = 8'hAA;
mem[16'h3938] = 8'hD5;
mem[16'h3939] = 8'hAA;
mem[16'h393A] = 8'hD5;
mem[16'h393B] = 8'hAA;
mem[16'h393C] = 8'hC5;
mem[16'h393D] = 8'hAA;
mem[16'h393E] = 8'hD5;
mem[16'h393F] = 8'hA8;
mem[16'h3940] = 8'hD5;
mem[16'h3941] = 8'h8A;
mem[16'h3942] = 8'hD5;
mem[16'h3943] = 8'hAA;
mem[16'h3944] = 8'hD5;
mem[16'h3945] = 8'hAA;
mem[16'h3946] = 8'hD5;
mem[16'h3947] = 8'hAA;
mem[16'h3948] = 8'hD5;
mem[16'h3949] = 8'hAA;
mem[16'h394A] = 8'hD5;
mem[16'h394B] = 8'hAA;
mem[16'h394C] = 8'h85;
mem[16'h394D] = 8'h00;
mem[16'h394E] = 8'h00;
mem[16'h394F] = 8'h2A;
mem[16'h3950] = 8'h00;
mem[16'h3951] = 8'hD8;
mem[16'h3952] = 8'h8D;
mem[16'h3953] = 8'h82;
mem[16'h3954] = 8'h00;
mem[16'h3955] = 8'h00;
mem[16'h3956] = 8'h00;
mem[16'h3957] = 8'h00;
mem[16'h3958] = 8'h00;
mem[16'h3959] = 8'h00;
mem[16'h395A] = 8'h00;
mem[16'h395B] = 8'hC0;
mem[16'h395C] = 8'hED;
mem[16'h395D] = 8'h90;
mem[16'h395E] = 8'h00;
mem[16'h395F] = 8'h00;
mem[16'h3960] = 8'h00;
mem[16'h3961] = 8'h00;
mem[16'h3962] = 8'h00;
mem[16'h3963] = 8'h00;
mem[16'h3964] = 8'h00;
mem[16'h3965] = 8'h00;
mem[16'h3966] = 8'hEC;
mem[16'h3967] = 8'h86;
mem[16'h3968] = 8'h81;
mem[16'h3969] = 8'h00;
mem[16'h396A] = 8'h00;
mem[16'h396B] = 8'h00;
mem[16'h396C] = 8'h00;
mem[16'h396D] = 8'h00;
mem[16'h396E] = 8'h00;
mem[16'h396F] = 8'h00;
mem[16'h3970] = 8'h00;
mem[16'h3971] = 8'h00;
mem[16'h3972] = 8'h00;
mem[16'h3973] = 8'h00;
mem[16'h3974] = 8'h00;
mem[16'h3975] = 8'h00;
mem[16'h3976] = 8'h00;
mem[16'h3977] = 8'h2A;
mem[16'h3978] = 8'h00;
mem[16'h3979] = 8'h00;
mem[16'h397A] = 8'h00;
mem[16'h397B] = 8'h00;
mem[16'h397C] = 8'h00;
mem[16'h397D] = 8'h00;
mem[16'h397E] = 8'h00;
mem[16'h397F] = 8'h00;
mem[16'h3980] = 8'hD5;
mem[16'h3981] = 8'hAA;
mem[16'h3982] = 8'hD5;
mem[16'h3983] = 8'hAA;
mem[16'h3984] = 8'hD5;
mem[16'h3985] = 8'hAA;
mem[16'h3986] = 8'hAD;
mem[16'h3987] = 8'hD5;
mem[16'h3988] = 8'hAA;
mem[16'h3989] = 8'hD5;
mem[16'h398A] = 8'hAA;
mem[16'h398B] = 8'hD5;
mem[16'h398C] = 8'hAA;
mem[16'h398D] = 8'hD5;
mem[16'h398E] = 8'hAA;
mem[16'h398F] = 8'hB5;
mem[16'h3990] = 8'hD5;
mem[16'h3991] = 8'hAA;
mem[16'h3992] = 8'hB5;
mem[16'h3993] = 8'hD5;
mem[16'h3994] = 8'hAA;
mem[16'h3995] = 8'hD5;
mem[16'h3996] = 8'hAA;
mem[16'h3997] = 8'hD5;
mem[16'h3998] = 8'hAA;
mem[16'h3999] = 8'hD5;
mem[16'h399A] = 8'hAA;
mem[16'h399B] = 8'hD5;
mem[16'h399C] = 8'hD5;
mem[16'h399D] = 8'hAA;
mem[16'h399E] = 8'hD5;
mem[16'h399F] = 8'hAA;
mem[16'h39A0] = 8'hD5;
mem[16'h39A1] = 8'hAA;
mem[16'h39A2] = 8'hD5;
mem[16'h39A3] = 8'hAA;
mem[16'h39A4] = 8'h85;
mem[16'h39A5] = 8'h00;
mem[16'h39A6] = 8'h00;
mem[16'h39A7] = 8'h00;
mem[16'h39A8] = 8'h0A;
mem[16'h39A9] = 8'h51;
mem[16'h39AA] = 8'h2A;
mem[16'h39AB] = 8'h10;
mem[16'h39AC] = 8'h28;
mem[16'h39AD] = 8'h45;
mem[16'h39AE] = 8'h2A;
mem[16'h39AF] = 8'h51;
mem[16'h39B0] = 8'h0A;
mem[16'h39B1] = 8'h51;
mem[16'h39B2] = 8'h2A;
mem[16'h39B3] = 8'h10;
mem[16'h39B4] = 8'h28;
mem[16'h39B5] = 8'h45;
mem[16'h39B6] = 8'h2A;
mem[16'h39B7] = 8'h51;
mem[16'h39B8] = 8'h0A;
mem[16'h39B9] = 8'h51;
mem[16'h39BA] = 8'h2A;
mem[16'h39BB] = 8'h10;
mem[16'h39BC] = 8'h28;
mem[16'h39BD] = 8'h45;
mem[16'h39BE] = 8'h2A;
mem[16'h39BF] = 8'h51;
mem[16'h39C0] = 8'h0A;
mem[16'h39C1] = 8'h51;
mem[16'h39C2] = 8'h2A;
mem[16'h39C3] = 8'h10;
mem[16'h39C4] = 8'h28;
mem[16'h39C5] = 8'h45;
mem[16'h39C6] = 8'h2A;
mem[16'h39C7] = 8'h51;
mem[16'h39C8] = 8'h0A;
mem[16'h39C9] = 8'h51;
mem[16'h39CA] = 8'h2A;
mem[16'h39CB] = 8'h10;
mem[16'h39CC] = 8'h08;
mem[16'h39CD] = 8'h00;
mem[16'h39CE] = 8'h00;
mem[16'h39CF] = 8'h2A;
mem[16'h39D0] = 8'h00;
mem[16'h39D1] = 8'h00;
mem[16'h39D2] = 8'h00;
mem[16'h39D3] = 8'h00;
mem[16'h39D4] = 8'h00;
mem[16'h39D5] = 8'h00;
mem[16'h39D6] = 8'h00;
mem[16'h39D7] = 8'h00;
mem[16'h39D8] = 8'h00;
mem[16'h39D9] = 8'h00;
mem[16'h39DA] = 8'h00;
mem[16'h39DB] = 8'h00;
mem[16'h39DC] = 8'h00;
mem[16'h39DD] = 8'h00;
mem[16'h39DE] = 8'h00;
mem[16'h39DF] = 8'h00;
mem[16'h39E0] = 8'h00;
mem[16'h39E1] = 8'h00;
mem[16'h39E2] = 8'h00;
mem[16'h39E3] = 8'h00;
mem[16'h39E4] = 8'h00;
mem[16'h39E5] = 8'h00;
mem[16'h39E6] = 8'h00;
mem[16'h39E7] = 8'h00;
mem[16'h39E8] = 8'h00;
mem[16'h39E9] = 8'h00;
mem[16'h39EA] = 8'h00;
mem[16'h39EB] = 8'h00;
mem[16'h39EC] = 8'h00;
mem[16'h39ED] = 8'h00;
mem[16'h39EE] = 8'h00;
mem[16'h39EF] = 8'h00;
mem[16'h39F0] = 8'h00;
mem[16'h39F1] = 8'h00;
mem[16'h39F2] = 8'h00;
mem[16'h39F3] = 8'h00;
mem[16'h39F4] = 8'h00;
mem[16'h39F5] = 8'h00;
mem[16'h39F6] = 8'h00;
mem[16'h39F7] = 8'h2A;
mem[16'h39F8] = 8'h00;
mem[16'h39F9] = 8'h00;
mem[16'h39FA] = 8'h00;
mem[16'h39FB] = 8'h00;
mem[16'h39FC] = 8'h00;
mem[16'h39FD] = 8'h00;
mem[16'h39FE] = 8'h00;
mem[16'h39FF] = 8'h00;
mem[16'h3A00] = 8'hD5;
mem[16'h3A01] = 8'hA8;
mem[16'h3A02] = 8'hD4;
mem[16'h3A03] = 8'h8A;
mem[16'h3A04] = 8'hC5;
mem[16'h3A05] = 8'hAA;
mem[16'h3A06] = 8'hD5;
mem[16'h3A07] = 8'hAA;
mem[16'h3A08] = 8'hD5;
mem[16'h3A09] = 8'hA2;
mem[16'h3A0A] = 8'hD1;
mem[16'h3A0B] = 8'hAA;
mem[16'h3A0C] = 8'h94;
mem[16'h3A0D] = 8'hAA;
mem[16'h3A0E] = 8'hD5;
mem[16'h3A0F] = 8'hAA;
mem[16'h3A10] = 8'hD5;
mem[16'h3A11] = 8'h8A;
mem[16'h3A12] = 8'hC5;
mem[16'h3A13] = 8'hAA;
mem[16'h3A14] = 8'hD1;
mem[16'h3A15] = 8'hA8;
mem[16'h3A16] = 8'hD5;
mem[16'h3A17] = 8'hAA;
mem[16'h3A18] = 8'hD5;
mem[16'h3A19] = 8'hAA;
mem[16'h3A1A] = 8'h94;
mem[16'h3A1B] = 8'hAA;
mem[16'h3A1C] = 8'hC5;
mem[16'h3A1D] = 8'hA2;
mem[16'h3A1E] = 8'hD5;
mem[16'h3A1F] = 8'hAA;
mem[16'h3A20] = 8'hD5;
mem[16'h3A21] = 8'hAA;
mem[16'h3A22] = 8'hD5;
mem[16'h3A23] = 8'hAA;
mem[16'h3A24] = 8'h85;
mem[16'h3A25] = 8'h00;
mem[16'h3A26] = 8'h7C;
mem[16'h3A27] = 8'h1F;
mem[16'h3A28] = 8'h0A;
mem[16'h3A29] = 8'h51;
mem[16'h3A2A] = 8'h2A;
mem[16'h3A2B] = 8'h10;
mem[16'h3A2C] = 8'h28;
mem[16'h3A2D] = 8'h45;
mem[16'h3A2E] = 8'h2A;
mem[16'h3A2F] = 8'h51;
mem[16'h3A30] = 8'h0A;
mem[16'h3A31] = 8'h51;
mem[16'h3A32] = 8'h2A;
mem[16'h3A33] = 8'h10;
mem[16'h3A34] = 8'h28;
mem[16'h3A35] = 8'h45;
mem[16'h3A36] = 8'h2A;
mem[16'h3A37] = 8'h51;
mem[16'h3A38] = 8'h0A;
mem[16'h3A39] = 8'h51;
mem[16'h3A3A] = 8'h2A;
mem[16'h3A3B] = 8'h10;
mem[16'h3A3C] = 8'h28;
mem[16'h3A3D] = 8'h45;
mem[16'h3A3E] = 8'h2A;
mem[16'h3A3F] = 8'h51;
mem[16'h3A40] = 8'h0A;
mem[16'h3A41] = 8'h51;
mem[16'h3A42] = 8'h2A;
mem[16'h3A43] = 8'h10;
mem[16'h3A44] = 8'h28;
mem[16'h3A45] = 8'h45;
mem[16'h3A46] = 8'h2A;
mem[16'h3A47] = 8'h51;
mem[16'h3A48] = 8'h0A;
mem[16'h3A49] = 8'h51;
mem[16'h3A4A] = 8'h2A;
mem[16'h3A4B] = 8'h10;
mem[16'h3A4C] = 8'h08;
mem[16'h3A4D] = 8'h00;
mem[16'h3A4E] = 8'h00;
mem[16'h3A4F] = 8'h2A;
mem[16'h3A50] = 8'h00;
mem[16'h3A51] = 8'h00;
mem[16'h3A52] = 8'h00;
mem[16'h3A53] = 8'h00;
mem[16'h3A54] = 8'h15;
mem[16'h3A55] = 8'h28;
mem[16'h3A56] = 8'h1D;
mem[16'h3A57] = 8'h00;
mem[16'h3A58] = 8'h00;
mem[16'h3A59] = 8'h00;
mem[16'h3A5A] = 8'h00;
mem[16'h3A5B] = 8'h00;
mem[16'h3A5C] = 8'h00;
mem[16'h3A5D] = 8'h00;
mem[16'h3A5E] = 8'h00;
mem[16'h3A5F] = 8'h00;
mem[16'h3A60] = 8'h00;
mem[16'h3A61] = 8'h00;
mem[16'h3A62] = 8'h15;
mem[16'h3A63] = 8'h28;
mem[16'h3A64] = 8'h1D;
mem[16'h3A65] = 8'h00;
mem[16'h3A66] = 8'h00;
mem[16'h3A67] = 8'h00;
mem[16'h3A68] = 8'h00;
mem[16'h3A69] = 8'h00;
mem[16'h3A6A] = 8'h00;
mem[16'h3A6B] = 8'h00;
mem[16'h3A6C] = 8'h00;
mem[16'h3A6D] = 8'h00;
mem[16'h3A6E] = 8'h00;
mem[16'h3A6F] = 8'h00;
mem[16'h3A70] = 8'h15;
mem[16'h3A71] = 8'h28;
mem[16'h3A72] = 8'h1D;
mem[16'h3A73] = 8'h00;
mem[16'h3A74] = 8'h00;
mem[16'h3A75] = 8'h00;
mem[16'h3A76] = 8'h00;
mem[16'h3A77] = 8'h2A;
mem[16'h3A78] = 8'h00;
mem[16'h3A79] = 8'h00;
mem[16'h3A7A] = 8'h00;
mem[16'h3A7B] = 8'h00;
mem[16'h3A7C] = 8'h00;
mem[16'h3A7D] = 8'h00;
mem[16'h3A7E] = 8'h00;
mem[16'h3A7F] = 8'h00;
mem[16'h3A80] = 8'hD5;
mem[16'h3A81] = 8'hA8;
mem[16'h3A82] = 8'hD4;
mem[16'h3A83] = 8'h8A;
mem[16'h3A84] = 8'hC5;
mem[16'h3A85] = 8'hAA;
mem[16'h3A86] = 8'hD5;
mem[16'h3A87] = 8'hAA;
mem[16'h3A88] = 8'hD5;
mem[16'h3A89] = 8'hA2;
mem[16'h3A8A] = 8'hD1;
mem[16'h3A8B] = 8'hAA;
mem[16'h3A8C] = 8'h94;
mem[16'h3A8D] = 8'hAA;
mem[16'h3A8E] = 8'hD5;
mem[16'h3A8F] = 8'hAA;
mem[16'h3A90] = 8'hD5;
mem[16'h3A91] = 8'h8A;
mem[16'h3A92] = 8'hC5;
mem[16'h3A93] = 8'hAA;
mem[16'h3A94] = 8'hD1;
mem[16'h3A95] = 8'hA8;
mem[16'h3A96] = 8'hD5;
mem[16'h3A97] = 8'hAA;
mem[16'h3A98] = 8'hD5;
mem[16'h3A99] = 8'hAA;
mem[16'h3A9A] = 8'h94;
mem[16'h3A9B] = 8'hAA;
mem[16'h3A9C] = 8'hC5;
mem[16'h3A9D] = 8'hA2;
mem[16'h3A9E] = 8'hD5;
mem[16'h3A9F] = 8'hAA;
mem[16'h3AA0] = 8'hD5;
mem[16'h3AA1] = 8'hAA;
mem[16'h3AA2] = 8'hD5;
mem[16'h3AA3] = 8'hAA;
mem[16'h3AA4] = 8'h85;
mem[16'h3AA5] = 8'h00;
mem[16'h3AA6] = 8'h60;
mem[16'h3AA7] = 8'h03;
mem[16'h3AA8] = 8'h00;
mem[16'h3AA9] = 8'h00;
mem[16'h3AAA] = 8'h1D;
mem[16'h3AAB] = 8'h55;
mem[16'h3AAC] = 8'h0A;
mem[16'h3AAD] = 8'h00;
mem[16'h3AAE] = 8'h00;
mem[16'h3AAF] = 8'h00;
mem[16'h3AB0] = 8'h00;
mem[16'h3AB1] = 8'h00;
mem[16'h3AB2] = 8'h00;
mem[16'h3AB3] = 8'h00;
mem[16'h3AB4] = 8'h00;
mem[16'h3AB5] = 8'h00;
mem[16'h3AB6] = 8'h00;
mem[16'h3AB7] = 8'h00;
mem[16'h3AB8] = 8'h1D;
mem[16'h3AB9] = 8'h55;
mem[16'h3ABA] = 8'h0A;
mem[16'h3ABB] = 8'h00;
mem[16'h3ABC] = 8'h00;
mem[16'h3ABD] = 8'h00;
mem[16'h3ABE] = 8'h00;
mem[16'h3ABF] = 8'h00;
mem[16'h3AC0] = 8'h00;
mem[16'h3AC1] = 8'h00;
mem[16'h3AC2] = 8'h00;
mem[16'h3AC3] = 8'h00;
mem[16'h3AC4] = 8'h00;
mem[16'h3AC5] = 8'h00;
mem[16'h3AC6] = 8'h00;
mem[16'h3AC7] = 8'h00;
mem[16'h3AC8] = 8'h00;
mem[16'h3AC9] = 8'h00;
mem[16'h3ACA] = 8'h00;
mem[16'h3ACB] = 8'h00;
mem[16'h3ACC] = 8'h00;
mem[16'h3ACD] = 8'h00;
mem[16'h3ACE] = 8'h00;
mem[16'h3ACF] = 8'h2A;
mem[16'h3AD0] = 8'h00;
mem[16'h3AD1] = 8'h00;
mem[16'h3AD2] = 8'h00;
mem[16'h3AD3] = 8'h00;
mem[16'h3AD4] = 8'h00;
mem[16'h3AD5] = 8'h00;
mem[16'h3AD6] = 8'h00;
mem[16'h3AD7] = 8'h00;
mem[16'h3AD8] = 8'h00;
mem[16'h3AD9] = 8'h00;
mem[16'h3ADA] = 8'h00;
mem[16'h3ADB] = 8'h00;
mem[16'h3ADC] = 8'h00;
mem[16'h3ADD] = 8'h00;
mem[16'h3ADE] = 8'h00;
mem[16'h3ADF] = 8'h00;
mem[16'h3AE0] = 8'h00;
mem[16'h3AE1] = 8'h00;
mem[16'h3AE2] = 8'h00;
mem[16'h3AE3] = 8'h00;
mem[16'h3AE4] = 8'h00;
mem[16'h3AE5] = 8'h00;
mem[16'h3AE6] = 8'h00;
mem[16'h3AE7] = 8'h00;
mem[16'h3AE8] = 8'h00;
mem[16'h3AE9] = 8'h00;
mem[16'h3AEA] = 8'h00;
mem[16'h3AEB] = 8'h00;
mem[16'h3AEC] = 8'h00;
mem[16'h3AED] = 8'h00;
mem[16'h3AEE] = 8'h00;
mem[16'h3AEF] = 8'h00;
mem[16'h3AF0] = 8'h00;
mem[16'h3AF1] = 8'h00;
mem[16'h3AF2] = 8'h00;
mem[16'h3AF3] = 8'h00;
mem[16'h3AF4] = 8'h00;
mem[16'h3AF5] = 8'h00;
mem[16'h3AF6] = 8'h00;
mem[16'h3AF7] = 8'h2A;
mem[16'h3AF8] = 8'h00;
mem[16'h3AF9] = 8'h00;
mem[16'h3AFA] = 8'h00;
mem[16'h3AFB] = 8'h00;
mem[16'h3AFC] = 8'h00;
mem[16'h3AFD] = 8'h00;
mem[16'h3AFE] = 8'h00;
mem[16'h3AFF] = 8'h00;
mem[16'h3B00] = 8'hAB;
mem[16'h3B01] = 8'hAD;
mem[16'h3B02] = 8'hD5;
mem[16'h3B03] = 8'hAA;
mem[16'h3B04] = 8'hD5;
mem[16'h3B05] = 8'hAA;
mem[16'h3B06] = 8'hD5;
mem[16'h3B07] = 8'hAA;
mem[16'h3B08] = 8'hD5;
mem[16'h3B09] = 8'hAA;
mem[16'h3B0A] = 8'hD5;
mem[16'h3B0B] = 8'hD5;
mem[16'h3B0C] = 8'hAA;
mem[16'h3B0D] = 8'hD5;
mem[16'h3B0E] = 8'hAA;
mem[16'h3B0F] = 8'hD5;
mem[16'h3B10] = 8'hAA;
mem[16'h3B11] = 8'hD5;
mem[16'h3B12] = 8'hAA;
mem[16'h3B13] = 8'hD5;
mem[16'h3B14] = 8'hAA;
mem[16'h3B15] = 8'hD5;
mem[16'h3B16] = 8'hAA;
mem[16'h3B17] = 8'hD5;
mem[16'h3B18] = 8'hAA;
mem[16'h3B19] = 8'hD5;
mem[16'h3B1A] = 8'hD5;
mem[16'h3B1B] = 8'hAA;
mem[16'h3B1C] = 8'hD5;
mem[16'h3B1D] = 8'hAA;
mem[16'h3B1E] = 8'hD5;
mem[16'h3B1F] = 8'hAA;
mem[16'h3B20] = 8'hD5;
mem[16'h3B21] = 8'hAA;
mem[16'h3B22] = 8'hD5;
mem[16'h3B23] = 8'hAA;
mem[16'h3B24] = 8'h85;
mem[16'h3B25] = 8'h00;
mem[16'h3B26] = 8'h44;
mem[16'h3B27] = 8'h12;
mem[16'h3B28] = 8'h00;
mem[16'h3B29] = 8'h00;
mem[16'h3B2A] = 8'h00;
mem[16'h3B2B] = 8'h00;
mem[16'h3B2C] = 8'h00;
mem[16'h3B2D] = 8'h00;
mem[16'h3B2E] = 8'h00;
mem[16'h3B2F] = 8'h00;
mem[16'h3B30] = 8'h00;
mem[16'h3B31] = 8'h00;
mem[16'h3B32] = 8'h00;
mem[16'h3B33] = 8'h00;
mem[16'h3B34] = 8'h00;
mem[16'h3B35] = 8'h00;
mem[16'h3B36] = 8'h00;
mem[16'h3B37] = 8'h00;
mem[16'h3B38] = 8'h00;
mem[16'h3B39] = 8'h00;
mem[16'h3B3A] = 8'h00;
mem[16'h3B3B] = 8'h00;
mem[16'h3B3C] = 8'h00;
mem[16'h3B3D] = 8'h00;
mem[16'h3B3E] = 8'h00;
mem[16'h3B3F] = 8'h00;
mem[16'h3B40] = 8'h00;
mem[16'h3B41] = 8'h00;
mem[16'h3B42] = 8'h00;
mem[16'h3B43] = 8'h00;
mem[16'h3B44] = 8'h00;
mem[16'h3B45] = 8'h00;
mem[16'h3B46] = 8'h00;
mem[16'h3B47] = 8'h00;
mem[16'h3B48] = 8'h00;
mem[16'h3B49] = 8'h00;
mem[16'h3B4A] = 8'h00;
mem[16'h3B4B] = 8'h00;
mem[16'h3B4C] = 8'h00;
mem[16'h3B4D] = 8'h00;
mem[16'h3B4E] = 8'h00;
mem[16'h3B4F] = 8'h2A;
mem[16'h3B50] = 8'h2A;
mem[16'h3B51] = 8'h45;
mem[16'h3B52] = 8'h2A;
mem[16'h3B53] = 8'h44;
mem[16'h3B54] = 8'h2A;
mem[16'h3B55] = 8'h41;
mem[16'h3B56] = 8'h20;
mem[16'h3B57] = 8'h15;
mem[16'h3B58] = 8'h2A;
mem[16'h3B59] = 8'h45;
mem[16'h3B5A] = 8'h2A;
mem[16'h3B5B] = 8'h44;
mem[16'h3B5C] = 8'h2A;
mem[16'h3B5D] = 8'h41;
mem[16'h3B5E] = 8'h20;
mem[16'h3B5F] = 8'h15;
mem[16'h3B60] = 8'h2A;
mem[16'h3B61] = 8'h45;
mem[16'h3B62] = 8'h74;
mem[16'h3B63] = 8'h17;
mem[16'h3B64] = 8'h2A;
mem[16'h3B65] = 8'h41;
mem[16'h3B66] = 8'h20;
mem[16'h3B67] = 8'h15;
mem[16'h3B68] = 8'h2A;
mem[16'h3B69] = 8'h45;
mem[16'h3B6A] = 8'h2A;
mem[16'h3B6B] = 8'h44;
mem[16'h3B6C] = 8'h2A;
mem[16'h3B6D] = 8'h41;
mem[16'h3B6E] = 8'h20;
mem[16'h3B6F] = 8'h15;
mem[16'h3B70] = 8'h2A;
mem[16'h3B71] = 8'h45;
mem[16'h3B72] = 8'h2A;
mem[16'h3B73] = 8'h44;
mem[16'h3B74] = 8'h0A;
mem[16'h3B75] = 8'h00;
mem[16'h3B76] = 8'h00;
mem[16'h3B77] = 8'h2A;
mem[16'h3B78] = 8'h00;
mem[16'h3B79] = 8'h00;
mem[16'h3B7A] = 8'h00;
mem[16'h3B7B] = 8'h00;
mem[16'h3B7C] = 8'h00;
mem[16'h3B7D] = 8'h00;
mem[16'h3B7E] = 8'h00;
mem[16'h3B7F] = 8'h00;
mem[16'h3B80] = 8'hD5;
mem[16'h3B81] = 8'hAA;
mem[16'h3B82] = 8'hD5;
mem[16'h3B83] = 8'hAA;
mem[16'h3B84] = 8'hD5;
mem[16'h3B85] = 8'hAA;
mem[16'h3B86] = 8'hD5;
mem[16'h3B87] = 8'hAA;
mem[16'h3B88] = 8'hD5;
mem[16'h3B89] = 8'hAA;
mem[16'h3B8A] = 8'hD5;
mem[16'h3B8B] = 8'hAA;
mem[16'h3B8C] = 8'hD5;
mem[16'h3B8D] = 8'hAA;
mem[16'h3B8E] = 8'hD5;
mem[16'h3B8F] = 8'hAA;
mem[16'h3B90] = 8'hD5;
mem[16'h3B91] = 8'hAA;
mem[16'h3B92] = 8'hD5;
mem[16'h3B93] = 8'hAA;
mem[16'h3B94] = 8'hD5;
mem[16'h3B95] = 8'hAA;
mem[16'h3B96] = 8'hD5;
mem[16'h3B97] = 8'hAA;
mem[16'h3B98] = 8'hD5;
mem[16'h3B99] = 8'hAA;
mem[16'h3B9A] = 8'hD5;
mem[16'h3B9B] = 8'hAA;
mem[16'h3B9C] = 8'hD5;
mem[16'h3B9D] = 8'hAA;
mem[16'h3B9E] = 8'hD5;
mem[16'h3B9F] = 8'hAA;
mem[16'h3BA0] = 8'hD5;
mem[16'h3BA1] = 8'hAA;
mem[16'h3BA2] = 8'hD5;
mem[16'h3BA3] = 8'hAA;
mem[16'h3BA4] = 8'h85;
mem[16'h3BA5] = 8'h00;
mem[16'h3BA6] = 8'h00;
mem[16'h3BA7] = 8'h00;
mem[16'h3BA8] = 8'h00;
mem[16'h3BA9] = 8'hB8;
mem[16'h3BAA] = 8'hD5;
mem[16'h3BAB] = 8'h82;
mem[16'h3BAC] = 8'h00;
mem[16'h3BAD] = 8'h00;
mem[16'h3BAE] = 8'h00;
mem[16'h3BAF] = 8'h00;
mem[16'h3BB0] = 8'h00;
mem[16'h3BB1] = 8'h00;
mem[16'h3BB2] = 8'h00;
mem[16'h3BB3] = 8'h00;
mem[16'h3BB4] = 8'h00;
mem[16'h3BB5] = 8'h00;
mem[16'h3BB6] = 8'h00;
mem[16'h3BB7] = 8'h00;
mem[16'h3BB8] = 8'h00;
mem[16'h3BB9] = 8'h00;
mem[16'h3BBA] = 8'h00;
mem[16'h3BBB] = 8'h00;
mem[16'h3BBC] = 8'h00;
mem[16'h3BBD] = 8'h00;
mem[16'h3BBE] = 8'h00;
mem[16'h3BBF] = 8'h00;
mem[16'h3BC0] = 8'h00;
mem[16'h3BC1] = 8'h00;
mem[16'h3BC2] = 8'h00;
mem[16'h3BC3] = 8'h00;
mem[16'h3BC4] = 8'h00;
mem[16'h3BC5] = 8'h00;
mem[16'h3BC6] = 8'h00;
mem[16'h3BC7] = 8'h00;
mem[16'h3BC8] = 8'h00;
mem[16'h3BC9] = 8'h00;
mem[16'h3BCA] = 8'h00;
mem[16'h3BCB] = 8'h00;
mem[16'h3BCC] = 8'h00;
mem[16'h3BCD] = 8'h00;
mem[16'h3BCE] = 8'h00;
mem[16'h3BCF] = 8'h2A;
mem[16'h3BD0] = 8'h00;
mem[16'h3BD1] = 8'h00;
mem[16'h3BD2] = 8'h00;
mem[16'h3BD3] = 8'h00;
mem[16'h3BD4] = 8'h00;
mem[16'h3BD5] = 8'h00;
mem[16'h3BD6] = 8'h00;
mem[16'h3BD7] = 8'h00;
mem[16'h3BD8] = 8'h00;
mem[16'h3BD9] = 8'h00;
mem[16'h3BDA] = 8'h00;
mem[16'h3BDB] = 8'h00;
mem[16'h3BDC] = 8'h00;
mem[16'h3BDD] = 8'h00;
mem[16'h3BDE] = 8'h00;
mem[16'h3BDF] = 8'h00;
mem[16'h3BE0] = 8'h00;
mem[16'h3BE1] = 8'h00;
mem[16'h3BE2] = 8'h00;
mem[16'h3BE3] = 8'h00;
mem[16'h3BE4] = 8'h00;
mem[16'h3BE5] = 8'h00;
mem[16'h3BE6] = 8'h00;
mem[16'h3BE7] = 8'h00;
mem[16'h3BE8] = 8'h00;
mem[16'h3BE9] = 8'h00;
mem[16'h3BEA] = 8'h00;
mem[16'h3BEB] = 8'h00;
mem[16'h3BEC] = 8'h00;
mem[16'h3BED] = 8'h00;
mem[16'h3BEE] = 8'h00;
mem[16'h3BEF] = 8'h00;
mem[16'h3BF0] = 8'h00;
mem[16'h3BF1] = 8'h00;
mem[16'h3BF2] = 8'h00;
mem[16'h3BF3] = 8'h00;
mem[16'h3BF4] = 8'h00;
mem[16'h3BF5] = 8'h42;
mem[16'h3BF6] = 8'h00;
mem[16'h3BF7] = 8'h00;
mem[16'h3BF8] = 8'h00;
mem[16'h3BF9] = 8'h00;
mem[16'h3BFA] = 8'h00;
mem[16'h3BFB] = 8'h00;
mem[16'h3BFC] = 8'h00;
mem[16'h3BFD] = 8'h00;
mem[16'h3BFE] = 8'h00;
mem[16'h3BFF] = 8'h00;
mem[16'h3C00] = 8'h00;
mem[16'h3C01] = 8'h00;
mem[16'h3C02] = 8'h00;
mem[16'h3C03] = 8'h00;
mem[16'h3C04] = 8'h00;
mem[16'h3C05] = 8'h00;
mem[16'h3C06] = 8'h00;
mem[16'h3C07] = 8'h00;
mem[16'h3C08] = 8'h00;
mem[16'h3C09] = 8'h00;
mem[16'h3C0A] = 8'h00;
mem[16'h3C0B] = 8'h00;
mem[16'h3C0C] = 8'h00;
mem[16'h3C0D] = 8'h00;
mem[16'h3C0E] = 8'h00;
mem[16'h3C0F] = 8'h00;
mem[16'h3C10] = 8'h00;
mem[16'h3C11] = 8'h00;
mem[16'h3C12] = 8'h00;
mem[16'h3C13] = 8'h00;
mem[16'h3C14] = 8'h00;
mem[16'h3C15] = 8'h00;
mem[16'h3C16] = 8'h00;
mem[16'h3C17] = 8'h00;
mem[16'h3C18] = 8'h00;
mem[16'h3C19] = 8'h00;
mem[16'h3C1A] = 8'h00;
mem[16'h3C1B] = 8'h00;
mem[16'h3C1C] = 8'h00;
mem[16'h3C1D] = 8'h00;
mem[16'h3C1E] = 8'h00;
mem[16'h3C1F] = 8'h00;
mem[16'h3C20] = 8'h00;
mem[16'h3C21] = 8'h00;
mem[16'h3C22] = 8'h00;
mem[16'h3C23] = 8'h00;
mem[16'h3C24] = 8'h00;
mem[16'h3C25] = 8'h00;
mem[16'h3C26] = 8'h60;
mem[16'h3C27] = 8'h03;
mem[16'h3C28] = 8'hD5;
mem[16'h3C29] = 8'hAA;
mem[16'h3C2A] = 8'hD5;
mem[16'h3C2B] = 8'hAA;
mem[16'h3C2C] = 8'hB5;
mem[16'h3C2D] = 8'hD5;
mem[16'h3C2E] = 8'hAA;
mem[16'h3C2F] = 8'hD5;
mem[16'h3C30] = 8'hAA;
mem[16'h3C31] = 8'hD5;
mem[16'h3C32] = 8'hAA;
mem[16'h3C33] = 8'hD5;
mem[16'h3C34] = 8'hD6;
mem[16'h3C35] = 8'hAA;
mem[16'h3C36] = 8'hD5;
mem[16'h3C37] = 8'hAA;
mem[16'h3C38] = 8'hD5;
mem[16'h3C39] = 8'hD5;
mem[16'h3C3A] = 8'hAA;
mem[16'h3C3B] = 8'hD5;
mem[16'h3C3C] = 8'hAA;
mem[16'h3C3D] = 8'hD5;
mem[16'h3C3E] = 8'hAA;
mem[16'h3C3F] = 8'hD5;
mem[16'h3C40] = 8'hDA;
mem[16'h3C41] = 8'hAA;
mem[16'h3C42] = 8'hD5;
mem[16'h3C43] = 8'hAA;
mem[16'h3C44] = 8'hAB;
mem[16'h3C45] = 8'hD5;
mem[16'h3C46] = 8'hAA;
mem[16'h3C47] = 8'hD5;
mem[16'h3C48] = 8'hAA;
mem[16'h3C49] = 8'hD5;
mem[16'h3C4A] = 8'hAA;
mem[16'h3C4B] = 8'hB5;
mem[16'h3C4C] = 8'h85;
mem[16'h3C4D] = 8'h00;
mem[16'h3C4E] = 8'h00;
mem[16'h3C4F] = 8'h2A;
mem[16'h3C50] = 8'h00;
mem[16'h3C51] = 8'h00;
mem[16'h3C52] = 8'h00;
mem[16'h3C53] = 8'h00;
mem[16'h3C54] = 8'h00;
mem[16'h3C55] = 8'h78;
mem[16'h3C56] = 8'h30;
mem[16'h3C57] = 8'h01;
mem[16'h3C58] = 8'h00;
mem[16'h3C59] = 8'h00;
mem[16'h3C5A] = 8'h00;
mem[16'h3C5B] = 8'h00;
mem[16'h3C5C] = 8'h00;
mem[16'h3C5D] = 8'h00;
mem[16'h3C5E] = 8'h00;
mem[16'h3C5F] = 8'h00;
mem[16'h3C60] = 8'h00;
mem[16'h3C61] = 8'h78;
mem[16'h3C62] = 8'h30;
mem[16'h3C63] = 8'h01;
mem[16'h3C64] = 8'h00;
mem[16'h3C65] = 8'h00;
mem[16'h3C66] = 8'h00;
mem[16'h3C67] = 8'h00;
mem[16'h3C68] = 8'h00;
mem[16'h3C69] = 8'h00;
mem[16'h3C6A] = 8'h00;
mem[16'h3C6B] = 8'h00;
mem[16'h3C6C] = 8'h00;
mem[16'h3C6D] = 8'h78;
mem[16'h3C6E] = 8'h30;
mem[16'h3C6F] = 8'h01;
mem[16'h3C70] = 8'h00;
mem[16'h3C71] = 8'h00;
mem[16'h3C72] = 8'h00;
mem[16'h3C73] = 8'h00;
mem[16'h3C74] = 8'h00;
mem[16'h3C75] = 8'h00;
mem[16'h3C76] = 8'h00;
mem[16'h3C77] = 8'h2A;
mem[16'h3C78] = 8'h00;
mem[16'h3C79] = 8'h00;
mem[16'h3C7A] = 8'h00;
mem[16'h3C7B] = 8'h00;
mem[16'h3C7C] = 8'h00;
mem[16'h3C7D] = 8'h00;
mem[16'h3C7E] = 8'h00;
mem[16'h3C7F] = 8'h00;
mem[16'h3C80] = 8'h28;
mem[16'h3C81] = 8'h15;
mem[16'h3C82] = 8'h08;
mem[16'h3C83] = 8'hAA;
mem[16'h3C84] = 8'hD5;
mem[16'h3C85] = 8'h55;
mem[16'h3C86] = 8'h28;
mem[16'h3C87] = 8'h45;
mem[16'h3C88] = 8'h28;
mem[16'h3C89] = 8'h15;
mem[16'h3C8A] = 8'hD5;
mem[16'h3C8B] = 8'hAA;
mem[16'h3C8C] = 8'h22;
mem[16'h3C8D] = 8'h55;
mem[16'h3C8E] = 8'h28;
mem[16'h3C8F] = 8'h45;
mem[16'h3C90] = 8'hD5;
mem[16'h3C91] = 8'hAA;
mem[16'h3C92] = 8'h08;
mem[16'h3C93] = 8'h54;
mem[16'h3C94] = 8'h22;
mem[16'h3C95] = 8'h55;
mem[16'h3C96] = 8'h28;
mem[16'h3C97] = 8'hAA;
mem[16'h3C98] = 8'hD5;
mem[16'h3C99] = 8'h15;
mem[16'h3C9A] = 8'h08;
mem[16'h3C9B] = 8'h54;
mem[16'h3C9C] = 8'h22;
mem[16'h3C9D] = 8'hAA;
mem[16'h3C9E] = 8'hD5;
mem[16'h3C9F] = 8'h45;
mem[16'h3CA0] = 8'h28;
mem[16'h3CA1] = 8'h15;
mem[16'h3CA2] = 8'h08;
mem[16'h3CA3] = 8'h54;
mem[16'h3CA4] = 8'h02;
mem[16'h3CA5] = 8'h00;
mem[16'h3CA6] = 8'h00;
mem[16'h3CA7] = 8'h00;
mem[16'h3CA8] = 8'hD5;
mem[16'h3CA9] = 8'hAA;
mem[16'h3CAA] = 8'hD5;
mem[16'h3CAB] = 8'hAA;
mem[16'h3CAC] = 8'hD5;
mem[16'h3CAD] = 8'hD6;
mem[16'h3CAE] = 8'hCA;
mem[16'h3CAF] = 8'hEA;
mem[16'h3CB0] = 8'hAA;
mem[16'h3CB1] = 8'hA9;
mem[16'h3CB2] = 8'hAD;
mem[16'h3CB3] = 8'h95;
mem[16'h3CB4] = 8'hD5;
mem[16'h3CB5] = 8'hAA;
mem[16'h3CB6] = 8'hD5;
mem[16'h3CB7] = 8'hAA;
mem[16'h3CB8] = 8'hD5;
mem[16'h3CB9] = 8'hAA;
mem[16'h3CBA] = 8'hD5;
mem[16'h3CBB] = 8'hAA;
mem[16'h3CBC] = 8'hAB;
mem[16'h3CBD] = 8'hA5;
mem[16'h3CBE] = 8'hB5;
mem[16'h3CBF] = 8'hD5;
mem[16'h3CC0] = 8'hD4;
mem[16'h3CC1] = 8'hD6;
mem[16'h3CC2] = 8'hCA;
mem[16'h3CC3] = 8'hAA;
mem[16'h3CC4] = 8'hD5;
mem[16'h3CC5] = 8'hAA;
mem[16'h3CC6] = 8'hD5;
mem[16'h3CC7] = 8'hAA;
mem[16'h3CC8] = 8'hD5;
mem[16'h3CC9] = 8'hAA;
mem[16'h3CCA] = 8'hD5;
mem[16'h3CCB] = 8'hAA;
mem[16'h3CCC] = 8'h85;
mem[16'h3CCD] = 8'h00;
mem[16'h3CCE] = 8'h00;
mem[16'h3CCF] = 8'h2A;
mem[16'h3CD0] = 8'h00;
mem[16'h3CD1] = 8'h00;
mem[16'h3CD2] = 8'h00;
mem[16'h3CD3] = 8'h00;
mem[16'h3CD4] = 8'h00;
mem[16'h3CD5] = 8'h00;
mem[16'h3CD6] = 8'h00;
mem[16'h3CD7] = 8'h00;
mem[16'h3CD8] = 8'h00;
mem[16'h3CD9] = 8'h00;
mem[16'h3CDA] = 8'h00;
mem[16'h3CDB] = 8'h00;
mem[16'h3CDC] = 8'h00;
mem[16'h3CDD] = 8'h00;
mem[16'h3CDE] = 8'h00;
mem[16'h3CDF] = 8'h00;
mem[16'h3CE0] = 8'h00;
mem[16'h3CE1] = 8'h00;
mem[16'h3CE2] = 8'h00;
mem[16'h3CE3] = 8'h00;
mem[16'h3CE4] = 8'h00;
mem[16'h3CE5] = 8'h00;
mem[16'h3CE6] = 8'h00;
mem[16'h3CE7] = 8'h00;
mem[16'h3CE8] = 8'h00;
mem[16'h3CE9] = 8'h00;
mem[16'h3CEA] = 8'h00;
mem[16'h3CEB] = 8'h00;
mem[16'h3CEC] = 8'h00;
mem[16'h3CED] = 8'h00;
mem[16'h3CEE] = 8'h00;
mem[16'h3CEF] = 8'h00;
mem[16'h3CF0] = 8'h00;
mem[16'h3CF1] = 8'h00;
mem[16'h3CF2] = 8'h00;
mem[16'h3CF3] = 8'h00;
mem[16'h3CF4] = 8'h00;
mem[16'h3CF5] = 8'h00;
mem[16'h3CF6] = 8'h00;
mem[16'h3CF7] = 8'h2A;
mem[16'h3CF8] = 8'h00;
mem[16'h3CF9] = 8'h00;
mem[16'h3CFA] = 8'h00;
mem[16'h3CFB] = 8'h00;
mem[16'h3CFC] = 8'h00;
mem[16'h3CFD] = 8'h00;
mem[16'h3CFE] = 8'h00;
mem[16'h3CFF] = 8'h00;
mem[16'h3D00] = 8'hD5;
mem[16'h3D01] = 8'hAA;
mem[16'h3D02] = 8'hD5;
mem[16'h3D03] = 8'hAA;
mem[16'h3D04] = 8'hD5;
mem[16'h3D05] = 8'hAA;
mem[16'h3D06] = 8'hB5;
mem[16'h3D07] = 8'hD5;
mem[16'h3D08] = 8'hAA;
mem[16'h3D09] = 8'hD5;
mem[16'h3D0A] = 8'hAA;
mem[16'h3D0B] = 8'hD5;
mem[16'h3D0C] = 8'hAA;
mem[16'h3D0D] = 8'hD5;
mem[16'h3D0E] = 8'hAA;
mem[16'h3D0F] = 8'hAD;
mem[16'h3D10] = 8'hD5;
mem[16'h3D11] = 8'hAA;
mem[16'h3D12] = 8'hD5;
mem[16'h3D13] = 8'hD5;
mem[16'h3D14] = 8'hAA;
mem[16'h3D15] = 8'hD5;
mem[16'h3D16] = 8'hAA;
mem[16'h3D17] = 8'hD5;
mem[16'h3D18] = 8'hAA;
mem[16'h3D19] = 8'hD5;
mem[16'h3D1A] = 8'hAA;
mem[16'h3D1B] = 8'hB5;
mem[16'h3D1C] = 8'hD5;
mem[16'h3D1D] = 8'hAA;
mem[16'h3D1E] = 8'hD5;
mem[16'h3D1F] = 8'hAA;
mem[16'h3D20] = 8'hD5;
mem[16'h3D21] = 8'hAA;
mem[16'h3D22] = 8'hD5;
mem[16'h3D23] = 8'hAA;
mem[16'h3D24] = 8'h85;
mem[16'h3D25] = 8'h00;
mem[16'h3D26] = 8'h74;
mem[16'h3D27] = 8'h17;
mem[16'h3D28] = 8'hD5;
mem[16'h3D29] = 8'hAA;
mem[16'h3D2A] = 8'hD5;
mem[16'h3D2B] = 8'hAA;
mem[16'h3D2C] = 8'hD5;
mem[16'h3D2D] = 8'hAA;
mem[16'h3D2E] = 8'hD5;
mem[16'h3D2F] = 8'hAA;
mem[16'h3D30] = 8'hD5;
mem[16'h3D31] = 8'hAA;
mem[16'h3D32] = 8'hD5;
mem[16'h3D33] = 8'hAA;
mem[16'h3D34] = 8'hD5;
mem[16'h3D35] = 8'hAA;
mem[16'h3D36] = 8'hD5;
mem[16'h3D37] = 8'hAA;
mem[16'h3D38] = 8'hD5;
mem[16'h3D39] = 8'hAA;
mem[16'h3D3A] = 8'hD5;
mem[16'h3D3B] = 8'hAA;
mem[16'h3D3C] = 8'hD5;
mem[16'h3D3D] = 8'hAA;
mem[16'h3D3E] = 8'hD5;
mem[16'h3D3F] = 8'hAA;
mem[16'h3D40] = 8'hD5;
mem[16'h3D41] = 8'hAA;
mem[16'h3D42] = 8'hD5;
mem[16'h3D43] = 8'hAA;
mem[16'h3D44] = 8'hD5;
mem[16'h3D45] = 8'hAA;
mem[16'h3D46] = 8'hD5;
mem[16'h3D47] = 8'hAA;
mem[16'h3D48] = 8'hD5;
mem[16'h3D49] = 8'hAA;
mem[16'h3D4A] = 8'hD5;
mem[16'h3D4B] = 8'hAA;
mem[16'h3D4C] = 8'h85;
mem[16'h3D4D] = 8'h00;
mem[16'h3D4E] = 8'h00;
mem[16'h3D4F] = 8'h2A;
mem[16'h3D50] = 8'h00;
mem[16'h3D51] = 8'hA8;
mem[16'h3D52] = 8'h95;
mem[16'h3D53] = 8'h81;
mem[16'h3D54] = 8'h00;
mem[16'h3D55] = 8'h00;
mem[16'h3D56] = 8'h00;
mem[16'h3D57] = 8'h00;
mem[16'h3D58] = 8'h00;
mem[16'h3D59] = 8'h00;
mem[16'h3D5A] = 8'h00;
mem[16'h3D5B] = 8'hC0;
mem[16'h3D5C] = 8'hAA;
mem[16'h3D5D] = 8'h89;
mem[16'h3D5E] = 8'h00;
mem[16'h3D5F] = 8'h00;
mem[16'h3D60] = 8'h00;
mem[16'h3D61] = 8'h00;
mem[16'h3D62] = 8'h00;
mem[16'h3D63] = 8'h00;
mem[16'h3D64] = 8'h00;
mem[16'h3D65] = 8'h00;
mem[16'h3D66] = 8'hD4;
mem[16'h3D67] = 8'hCA;
mem[16'h3D68] = 8'h80;
mem[16'h3D69] = 8'h00;
mem[16'h3D6A] = 8'h00;
mem[16'h3D6B] = 8'h00;
mem[16'h3D6C] = 8'h00;
mem[16'h3D6D] = 8'h00;
mem[16'h3D6E] = 8'h00;
mem[16'h3D6F] = 8'h00;
mem[16'h3D70] = 8'h00;
mem[16'h3D71] = 8'h00;
mem[16'h3D72] = 8'h00;
mem[16'h3D73] = 8'h00;
mem[16'h3D74] = 8'h00;
mem[16'h3D75] = 8'h00;
mem[16'h3D76] = 8'h00;
mem[16'h3D77] = 8'h2A;
mem[16'h3D78] = 8'h00;
mem[16'h3D79] = 8'h00;
mem[16'h3D7A] = 8'h00;
mem[16'h3D7B] = 8'h00;
mem[16'h3D7C] = 8'h00;
mem[16'h3D7D] = 8'h00;
mem[16'h3D7E] = 8'h00;
mem[16'h3D7F] = 8'h00;
mem[16'h3D80] = 8'hD5;
mem[16'h3D81] = 8'hAA;
mem[16'h3D82] = 8'hD5;
mem[16'h3D83] = 8'hAA;
mem[16'h3D84] = 8'hD5;
mem[16'h3D85] = 8'hAA;
mem[16'h3D86] = 8'hB5;
mem[16'h3D87] = 8'hD5;
mem[16'h3D88] = 8'hAA;
mem[16'h3D89] = 8'hD5;
mem[16'h3D8A] = 8'hAA;
mem[16'h3D8B] = 8'hD5;
mem[16'h3D8C] = 8'hAA;
mem[16'h3D8D] = 8'hD5;
mem[16'h3D8E] = 8'hAA;
mem[16'h3D8F] = 8'hAD;
mem[16'h3D90] = 8'hD5;
mem[16'h3D91] = 8'hAA;
mem[16'h3D92] = 8'hD5;
mem[16'h3D93] = 8'hD5;
mem[16'h3D94] = 8'hAA;
mem[16'h3D95] = 8'hD5;
mem[16'h3D96] = 8'hAA;
mem[16'h3D97] = 8'hD5;
mem[16'h3D98] = 8'hAA;
mem[16'h3D99] = 8'hD5;
mem[16'h3D9A] = 8'hAA;
mem[16'h3D9B] = 8'hB5;
mem[16'h3D9C] = 8'hD5;
mem[16'h3D9D] = 8'hAA;
mem[16'h3D9E] = 8'hD5;
mem[16'h3D9F] = 8'hAA;
mem[16'h3DA0] = 8'hD5;
mem[16'h3DA1] = 8'hAA;
mem[16'h3DA2] = 8'hD5;
mem[16'h3DA3] = 8'hAA;
mem[16'h3DA4] = 8'h85;
mem[16'h3DA5] = 8'h00;
mem[16'h3DA6] = 8'h40;
mem[16'h3DA7] = 8'h01;
mem[16'h3DA8] = 8'h0A;
mem[16'h3DA9] = 8'h04;
mem[16'h3DAA] = 8'h2A;
mem[16'h3DAB] = 8'h51;
mem[16'h3DAC] = 8'h2A;
mem[16'h3DAD] = 8'h54;
mem[16'h3DAE] = 8'h22;
mem[16'h3DAF] = 8'h54;
mem[16'h3DB0] = 8'h0A;
mem[16'h3DB1] = 8'h04;
mem[16'h3DB2] = 8'h2A;
mem[16'h3DB3] = 8'h51;
mem[16'h3DB4] = 8'h2A;
mem[16'h3DB5] = 8'h54;
mem[16'h3DB6] = 8'h22;
mem[16'h3DB7] = 8'h54;
mem[16'h3DB8] = 8'h0A;
mem[16'h3DB9] = 8'h04;
mem[16'h3DBA] = 8'h2A;
mem[16'h3DBB] = 8'h51;
mem[16'h3DBC] = 8'h2A;
mem[16'h3DBD] = 8'h54;
mem[16'h3DBE] = 8'h22;
mem[16'h3DBF] = 8'h54;
mem[16'h3DC0] = 8'h0A;
mem[16'h3DC1] = 8'h04;
mem[16'h3DC2] = 8'h2A;
mem[16'h3DC3] = 8'h51;
mem[16'h3DC4] = 8'h2A;
mem[16'h3DC5] = 8'h54;
mem[16'h3DC6] = 8'h22;
mem[16'h3DC7] = 8'h54;
mem[16'h3DC8] = 8'h0A;
mem[16'h3DC9] = 8'h04;
mem[16'h3DCA] = 8'h2A;
mem[16'h3DCB] = 8'h51;
mem[16'h3DCC] = 8'h0A;
mem[16'h3DCD] = 8'h00;
mem[16'h3DCE] = 8'h00;
mem[16'h3DCF] = 8'h2A;
mem[16'h3DD0] = 8'h00;
mem[16'h3DD1] = 8'h00;
mem[16'h3DD2] = 8'h00;
mem[16'h3DD3] = 8'h00;
mem[16'h3DD4] = 8'h00;
mem[16'h3DD5] = 8'h00;
mem[16'h3DD6] = 8'h00;
mem[16'h3DD7] = 8'h00;
mem[16'h3DD8] = 8'h00;
mem[16'h3DD9] = 8'h00;
mem[16'h3DDA] = 8'h00;
mem[16'h3DDB] = 8'h00;
mem[16'h3DDC] = 8'h00;
mem[16'h3DDD] = 8'h00;
mem[16'h3DDE] = 8'h00;
mem[16'h3DDF] = 8'h00;
mem[16'h3DE0] = 8'h00;
mem[16'h3DE1] = 8'h00;
mem[16'h3DE2] = 8'h00;
mem[16'h3DE3] = 8'h00;
mem[16'h3DE4] = 8'h00;
mem[16'h3DE5] = 8'h00;
mem[16'h3DE6] = 8'h00;
mem[16'h3DE7] = 8'h00;
mem[16'h3DE8] = 8'h00;
mem[16'h3DE9] = 8'h00;
mem[16'h3DEA] = 8'h00;
mem[16'h3DEB] = 8'h00;
mem[16'h3DEC] = 8'h00;
mem[16'h3DED] = 8'h00;
mem[16'h3DEE] = 8'h00;
mem[16'h3DEF] = 8'h00;
mem[16'h3DF0] = 8'h00;
mem[16'h3DF1] = 8'h00;
mem[16'h3DF2] = 8'h00;
mem[16'h3DF3] = 8'h00;
mem[16'h3DF4] = 8'h00;
mem[16'h3DF5] = 8'h00;
mem[16'h3DF6] = 8'h00;
mem[16'h3DF7] = 8'h2A;
mem[16'h3DF8] = 8'h00;
mem[16'h3DF9] = 8'h00;
mem[16'h3DFA] = 8'h00;
mem[16'h3DFB] = 8'h00;
mem[16'h3DFC] = 8'h00;
mem[16'h3DFD] = 8'h00;
mem[16'h3DFE] = 8'h00;
mem[16'h3DFF] = 8'h00;
mem[16'h3E00] = 8'hD5;
mem[16'h3E01] = 8'h94;
mem[16'h3E02] = 8'hD4;
mem[16'h3E03] = 8'hCA;
mem[16'h3E04] = 8'hC2;
mem[16'h3E05] = 8'hAA;
mem[16'h3E06] = 8'hD5;
mem[16'h3E07] = 8'hAA;
mem[16'h3E08] = 8'hD5;
mem[16'h3E09] = 8'hD2;
mem[16'h3E0A] = 8'hD0;
mem[16'h3E0B] = 8'hAA;
mem[16'h3E0C] = 8'h8A;
mem[16'h3E0D] = 8'hAA;
mem[16'h3E0E] = 8'hD5;
mem[16'h3E0F] = 8'hAA;
mem[16'h3E10] = 8'hD5;
mem[16'h3E11] = 8'hCA;
mem[16'h3E12] = 8'hC2;
mem[16'h3E13] = 8'hAA;
mem[16'h3E14] = 8'hA9;
mem[16'h3E15] = 8'hA8;
mem[16'h3E16] = 8'hD5;
mem[16'h3E17] = 8'hAA;
mem[16'h3E18] = 8'hD5;
mem[16'h3E19] = 8'hAA;
mem[16'h3E1A] = 8'h8A;
mem[16'h3E1B] = 8'hAA;
mem[16'h3E1C] = 8'hA5;
mem[16'h3E1D] = 8'hA1;
mem[16'h3E1E] = 8'hD5;
mem[16'h3E1F] = 8'hAA;
mem[16'h3E20] = 8'hD5;
mem[16'h3E21] = 8'hAA;
mem[16'h3E22] = 8'hD5;
mem[16'h3E23] = 8'hAA;
mem[16'h3E24] = 8'h85;
mem[16'h3E25] = 8'h00;
mem[16'h3E26] = 8'h7C;
mem[16'h3E27] = 8'h1F;
mem[16'h3E28] = 8'h2A;
mem[16'h3E29] = 8'h54;
mem[16'h3E2A] = 8'h0A;
mem[16'h3E2B] = 8'h55;
mem[16'h3E2C] = 8'h08;
mem[16'h3E2D] = 8'h55;
mem[16'h3E2E] = 8'h02;
mem[16'h3E2F] = 8'h41;
mem[16'h3E30] = 8'h2A;
mem[16'h3E31] = 8'h54;
mem[16'h3E32] = 8'h0A;
mem[16'h3E33] = 8'h55;
mem[16'h3E34] = 8'h08;
mem[16'h3E35] = 8'h55;
mem[16'h3E36] = 8'h02;
mem[16'h3E37] = 8'h41;
mem[16'h3E38] = 8'h2A;
mem[16'h3E39] = 8'h54;
mem[16'h3E3A] = 8'h0A;
mem[16'h3E3B] = 8'h55;
mem[16'h3E3C] = 8'h08;
mem[16'h3E3D] = 8'h55;
mem[16'h3E3E] = 8'h02;
mem[16'h3E3F] = 8'h41;
mem[16'h3E40] = 8'h2A;
mem[16'h3E41] = 8'h54;
mem[16'h3E42] = 8'h0A;
mem[16'h3E43] = 8'h55;
mem[16'h3E44] = 8'h08;
mem[16'h3E45] = 8'h55;
mem[16'h3E46] = 8'h02;
mem[16'h3E47] = 8'h41;
mem[16'h3E48] = 8'h2A;
mem[16'h3E49] = 8'h54;
mem[16'h3E4A] = 8'h0A;
mem[16'h3E4B] = 8'h55;
mem[16'h3E4C] = 8'h08;
mem[16'h3E4D] = 8'h00;
mem[16'h3E4E] = 8'h00;
mem[16'h3E4F] = 8'h2A;
mem[16'h3E50] = 8'h00;
mem[16'h3E51] = 8'h00;
mem[16'h3E52] = 8'h00;
mem[16'h3E53] = 8'h00;
mem[16'h3E54] = 8'h15;
mem[16'h3E55] = 8'h28;
mem[16'h3E56] = 8'h01;
mem[16'h3E57] = 8'h00;
mem[16'h3E58] = 8'h00;
mem[16'h3E59] = 8'h00;
mem[16'h3E5A] = 8'h00;
mem[16'h3E5B] = 8'h00;
mem[16'h3E5C] = 8'h00;
mem[16'h3E5D] = 8'h00;
mem[16'h3E5E] = 8'h00;
mem[16'h3E5F] = 8'h00;
mem[16'h3E60] = 8'h00;
mem[16'h3E61] = 8'h00;
mem[16'h3E62] = 8'h15;
mem[16'h3E63] = 8'h28;
mem[16'h3E64] = 8'h01;
mem[16'h3E65] = 8'h00;
mem[16'h3E66] = 8'h00;
mem[16'h3E67] = 8'h00;
mem[16'h3E68] = 8'h00;
mem[16'h3E69] = 8'h00;
mem[16'h3E6A] = 8'h00;
mem[16'h3E6B] = 8'h00;
mem[16'h3E6C] = 8'h00;
mem[16'h3E6D] = 8'h00;
mem[16'h3E6E] = 8'h00;
mem[16'h3E6F] = 8'h00;
mem[16'h3E70] = 8'h15;
mem[16'h3E71] = 8'h28;
mem[16'h3E72] = 8'h01;
mem[16'h3E73] = 8'h00;
mem[16'h3E74] = 8'h00;
mem[16'h3E75] = 8'h00;
mem[16'h3E76] = 8'h00;
mem[16'h3E77] = 8'h2A;
mem[16'h3E78] = 8'h00;
mem[16'h3E79] = 8'h00;
mem[16'h3E7A] = 8'h00;
mem[16'h3E7B] = 8'h00;
mem[16'h3E7C] = 8'h00;
mem[16'h3E7D] = 8'h00;
mem[16'h3E7E] = 8'h00;
mem[16'h3E7F] = 8'h00;
mem[16'h3E80] = 8'hD5;
mem[16'h3E81] = 8'hA8;
mem[16'h3E82] = 8'hD5;
mem[16'h3E83] = 8'h8A;
mem[16'h3E84] = 8'hD5;
mem[16'h3E85] = 8'hAA;
mem[16'h3E86] = 8'hD5;
mem[16'h3E87] = 8'hAA;
mem[16'h3E88] = 8'hD5;
mem[16'h3E89] = 8'hA2;
mem[16'h3E8A] = 8'hD5;
mem[16'h3E8B] = 8'hAA;
mem[16'h3E8C] = 8'hD4;
mem[16'h3E8D] = 8'hAA;
mem[16'h3E8E] = 8'hD5;
mem[16'h3E8F] = 8'hAA;
mem[16'h3E90] = 8'hD5;
mem[16'h3E91] = 8'h8A;
mem[16'h3E92] = 8'hD5;
mem[16'h3E93] = 8'hAA;
mem[16'h3E94] = 8'hD1;
mem[16'h3E95] = 8'hAA;
mem[16'h3E96] = 8'hD5;
mem[16'h3E97] = 8'hAA;
mem[16'h3E98] = 8'hD5;
mem[16'h3E99] = 8'hAA;
mem[16'h3E9A] = 8'hD4;
mem[16'h3E9B] = 8'hAA;
mem[16'h3E9C] = 8'hC5;
mem[16'h3E9D] = 8'hAA;
mem[16'h3E9E] = 8'hD5;
mem[16'h3E9F] = 8'hAA;
mem[16'h3EA0] = 8'hD5;
mem[16'h3EA1] = 8'hAA;
mem[16'h3EA2] = 8'hD5;
mem[16'h3EA3] = 8'hAA;
mem[16'h3EA4] = 8'h85;
mem[16'h3EA5] = 8'h00;
mem[16'h3EA6] = 8'h60;
mem[16'h3EA7] = 8'h03;
mem[16'h3EA8] = 8'h00;
mem[16'h3EA9] = 8'h00;
mem[16'h3EAA] = 8'h7D;
mem[16'h3EAB] = 8'h55;
mem[16'h3EAC] = 8'h0A;
mem[16'h3EAD] = 8'h00;
mem[16'h3EAE] = 8'h00;
mem[16'h3EAF] = 8'h00;
mem[16'h3EB0] = 8'h00;
mem[16'h3EB1] = 8'h00;
mem[16'h3EB2] = 8'h00;
mem[16'h3EB3] = 8'h00;
mem[16'h3EB4] = 8'h00;
mem[16'h3EB5] = 8'h00;
mem[16'h3EB6] = 8'h00;
mem[16'h3EB7] = 8'h00;
mem[16'h3EB8] = 8'h7D;
mem[16'h3EB9] = 8'h55;
mem[16'h3EBA] = 8'h0A;
mem[16'h3EBB] = 8'h00;
mem[16'h3EBC] = 8'h00;
mem[16'h3EBD] = 8'h00;
mem[16'h3EBE] = 8'h00;
mem[16'h3EBF] = 8'h00;
mem[16'h3EC0] = 8'h00;
mem[16'h3EC1] = 8'h00;
mem[16'h3EC2] = 8'h00;
mem[16'h3EC3] = 8'h00;
mem[16'h3EC4] = 8'h00;
mem[16'h3EC5] = 8'h00;
mem[16'h3EC6] = 8'h00;
mem[16'h3EC7] = 8'h00;
mem[16'h3EC8] = 8'h00;
mem[16'h3EC9] = 8'h00;
mem[16'h3ECA] = 8'h00;
mem[16'h3ECB] = 8'h00;
mem[16'h3ECC] = 8'h00;
mem[16'h3ECD] = 8'h00;
mem[16'h3ECE] = 8'h00;
mem[16'h3ECF] = 8'h2A;
mem[16'h3ED0] = 8'h0A;
mem[16'h3ED1] = 8'h51;
mem[16'h3ED2] = 8'h2A;
mem[16'h3ED3] = 8'h10;
mem[16'h3ED4] = 8'h28;
mem[16'h3ED5] = 8'h45;
mem[16'h3ED6] = 8'h2A;
mem[16'h3ED7] = 8'h51;
mem[16'h3ED8] = 8'h0A;
mem[16'h3ED9] = 8'h51;
mem[16'h3EDA] = 8'h2A;
mem[16'h3EDB] = 8'h10;
mem[16'h3EDC] = 8'h28;
mem[16'h3EDD] = 8'h45;
mem[16'h3EDE] = 8'h2A;
mem[16'h3EDF] = 8'h51;
mem[16'h3EE0] = 8'h0A;
mem[16'h3EE1] = 8'h51;
mem[16'h3EE2] = 8'h00;
mem[16'h3EE3] = 8'h00;
mem[16'h3EE4] = 8'h28;
mem[16'h3EE5] = 8'h45;
mem[16'h3EE6] = 8'h2A;
mem[16'h3EE7] = 8'h51;
mem[16'h3EE8] = 8'h0A;
mem[16'h3EE9] = 8'h51;
mem[16'h3EEA] = 8'h2A;
mem[16'h3EEB] = 8'h10;
mem[16'h3EEC] = 8'h28;
mem[16'h3EED] = 8'h45;
mem[16'h3EEE] = 8'h2A;
mem[16'h3EEF] = 8'h51;
mem[16'h3EF0] = 8'h0A;
mem[16'h3EF1] = 8'h51;
mem[16'h3EF2] = 8'h2A;
mem[16'h3EF3] = 8'h10;
mem[16'h3EF4] = 8'h08;
mem[16'h3EF5] = 8'h00;
mem[16'h3EF6] = 8'h00;
mem[16'h3EF7] = 8'h2A;
mem[16'h3EF8] = 8'h00;
mem[16'h3EF9] = 8'h00;
mem[16'h3EFA] = 8'h00;
mem[16'h3EFB] = 8'h00;
mem[16'h3EFC] = 8'h00;
mem[16'h3EFD] = 8'h00;
mem[16'h3EFE] = 8'h00;
mem[16'h3EFF] = 8'h00;
mem[16'h3F00] = 8'hAB;
mem[16'h3F01] = 8'hAD;
mem[16'h3F02] = 8'hD5;
mem[16'h3F03] = 8'hAA;
mem[16'h3F04] = 8'hD5;
mem[16'h3F05] = 8'hAA;
mem[16'h3F06] = 8'hD5;
mem[16'h3F07] = 8'hAA;
mem[16'h3F08] = 8'hD5;
mem[16'h3F09] = 8'hAA;
mem[16'h3F0A] = 8'hD5;
mem[16'h3F0B] = 8'hD5;
mem[16'h3F0C] = 8'hAA;
mem[16'h3F0D] = 8'hD5;
mem[16'h3F0E] = 8'hAA;
mem[16'h3F0F] = 8'hD5;
mem[16'h3F10] = 8'hAA;
mem[16'h3F11] = 8'hD5;
mem[16'h3F12] = 8'hAA;
mem[16'h3F13] = 8'hD5;
mem[16'h3F14] = 8'hAA;
mem[16'h3F15] = 8'hD5;
mem[16'h3F16] = 8'hAA;
mem[16'h3F17] = 8'hD5;
mem[16'h3F18] = 8'hAA;
mem[16'h3F19] = 8'hD5;
mem[16'h3F1A] = 8'hD5;
mem[16'h3F1B] = 8'hAA;
mem[16'h3F1C] = 8'hD5;
mem[16'h3F1D] = 8'hAA;
mem[16'h3F1E] = 8'hD5;
mem[16'h3F1F] = 8'hAA;
mem[16'h3F20] = 8'hD5;
mem[16'h3F21] = 8'hAA;
mem[16'h3F22] = 8'hD5;
mem[16'h3F23] = 8'hAA;
mem[16'h3F24] = 8'h85;
mem[16'h3F25] = 8'h00;
mem[16'h3F26] = 8'h0E;
mem[16'h3F27] = 8'h38;
mem[16'h3F28] = 8'h00;
mem[16'h3F29] = 8'h00;
mem[16'h3F2A] = 8'h00;
mem[16'h3F2B] = 8'h00;
mem[16'h3F2C] = 8'h00;
mem[16'h3F2D] = 8'h00;
mem[16'h3F2E] = 8'h00;
mem[16'h3F2F] = 8'h00;
mem[16'h3F30] = 8'h00;
mem[16'h3F31] = 8'h00;
mem[16'h3F32] = 8'h00;
mem[16'h3F33] = 8'h00;
mem[16'h3F34] = 8'h00;
mem[16'h3F35] = 8'h00;
mem[16'h3F36] = 8'h00;
mem[16'h3F37] = 8'h00;
mem[16'h3F38] = 8'h00;
mem[16'h3F39] = 8'h00;
mem[16'h3F3A] = 8'h00;
mem[16'h3F3B] = 8'h00;
mem[16'h3F3C] = 8'h00;
mem[16'h3F3D] = 8'h00;
mem[16'h3F3E] = 8'h00;
mem[16'h3F3F] = 8'h00;
mem[16'h3F40] = 8'h00;
mem[16'h3F41] = 8'h00;
mem[16'h3F42] = 8'h00;
mem[16'h3F43] = 8'h00;
mem[16'h3F44] = 8'h00;
mem[16'h3F45] = 8'h00;
mem[16'h3F46] = 8'h00;
mem[16'h3F47] = 8'h00;
mem[16'h3F48] = 8'h00;
mem[16'h3F49] = 8'h00;
mem[16'h3F4A] = 8'h00;
mem[16'h3F4B] = 8'h00;
mem[16'h3F4C] = 8'h00;
mem[16'h3F4D] = 8'h00;
mem[16'h3F4E] = 8'h00;
mem[16'h3F4F] = 8'h2A;
mem[16'h3F50] = 8'h0A;
mem[16'h3F51] = 8'h04;
mem[16'h3F52] = 8'h2A;
mem[16'h3F53] = 8'h51;
mem[16'h3F54] = 8'h2A;
mem[16'h3F55] = 8'h54;
mem[16'h3F56] = 8'h22;
mem[16'h3F57] = 8'h54;
mem[16'h3F58] = 8'h0A;
mem[16'h3F59] = 8'h04;
mem[16'h3F5A] = 8'h2A;
mem[16'h3F5B] = 8'h51;
mem[16'h3F5C] = 8'h2A;
mem[16'h3F5D] = 8'h54;
mem[16'h3F5E] = 8'h22;
mem[16'h3F5F] = 8'h54;
mem[16'h3F60] = 8'h0A;
mem[16'h3F61] = 8'h04;
mem[16'h3F62] = 8'h7C;
mem[16'h3F63] = 8'h1F;
mem[16'h3F64] = 8'h2A;
mem[16'h3F65] = 8'h54;
mem[16'h3F66] = 8'h22;
mem[16'h3F67] = 8'h54;
mem[16'h3F68] = 8'h0A;
mem[16'h3F69] = 8'h04;
mem[16'h3F6A] = 8'h2A;
mem[16'h3F6B] = 8'h51;
mem[16'h3F6C] = 8'h2A;
mem[16'h3F6D] = 8'h54;
mem[16'h3F6E] = 8'h22;
mem[16'h3F6F] = 8'h54;
mem[16'h3F70] = 8'h0A;
mem[16'h3F71] = 8'h04;
mem[16'h3F72] = 8'h2A;
mem[16'h3F73] = 8'h51;
mem[16'h3F74] = 8'h0A;
mem[16'h3F75] = 8'h00;
mem[16'h3F76] = 8'h00;
mem[16'h3F77] = 8'h2A;
mem[16'h3F78] = 8'h00;
mem[16'h3F79] = 8'h00;
mem[16'h3F7A] = 8'h00;
mem[16'h3F7B] = 8'h00;
mem[16'h3F7C] = 8'h00;
mem[16'h3F7D] = 8'h00;
mem[16'h3F7E] = 8'h00;
mem[16'h3F7F] = 8'h00;
mem[16'h3F80] = 8'hD5;
mem[16'h3F81] = 8'hAA;
mem[16'h3F82] = 8'hD5;
mem[16'h3F83] = 8'hAA;
mem[16'h3F84] = 8'hD5;
mem[16'h3F85] = 8'hAA;
mem[16'h3F86] = 8'hD5;
mem[16'h3F87] = 8'hAA;
mem[16'h3F88] = 8'hD5;
mem[16'h3F89] = 8'hAA;
mem[16'h3F8A] = 8'hD5;
mem[16'h3F8B] = 8'hAA;
mem[16'h3F8C] = 8'hD5;
mem[16'h3F8D] = 8'hAA;
mem[16'h3F8E] = 8'hD5;
mem[16'h3F8F] = 8'hAA;
mem[16'h3F90] = 8'hD5;
mem[16'h3F91] = 8'hAA;
mem[16'h3F92] = 8'hD5;
mem[16'h3F93] = 8'hAA;
mem[16'h3F94] = 8'hD5;
mem[16'h3F95] = 8'hAA;
mem[16'h3F96] = 8'hD5;
mem[16'h3F97] = 8'hAA;
mem[16'h3F98] = 8'hD5;
mem[16'h3F99] = 8'hAA;
mem[16'h3F9A] = 8'hD5;
mem[16'h3F9B] = 8'hAA;
mem[16'h3F9C] = 8'hD5;
mem[16'h3F9D] = 8'hAA;
mem[16'h3F9E] = 8'hD5;
mem[16'h3F9F] = 8'hAA;
mem[16'h3FA0] = 8'hD5;
mem[16'h3FA1] = 8'hAA;
mem[16'h3FA2] = 8'hD5;
mem[16'h3FA3] = 8'hAA;
mem[16'h3FA4] = 8'h85;
mem[16'h3FA5] = 8'h00;
mem[16'h3FA6] = 8'h00;
mem[16'h3FA7] = 8'h00;
mem[16'h3FA8] = 8'h00;
mem[16'h3FA9] = 8'hA0;
mem[16'h3FAA] = 8'h94;
mem[16'h3FAB] = 8'h81;
mem[16'h3FAC] = 8'h00;
mem[16'h3FAD] = 8'h00;
mem[16'h3FAE] = 8'h00;
mem[16'h3FAF] = 8'h00;
mem[16'h3FB0] = 8'h00;
mem[16'h3FB1] = 8'h00;
mem[16'h3FB2] = 8'h00;
mem[16'h3FB3] = 8'h00;
mem[16'h3FB4] = 8'h00;
mem[16'h3FB5] = 8'h00;
mem[16'h3FB6] = 8'h00;
mem[16'h3FB7] = 8'h00;
mem[16'h3FB8] = 8'h00;
mem[16'h3FB9] = 8'h00;
mem[16'h3FBA] = 8'h00;
mem[16'h3FBB] = 8'h00;
mem[16'h3FBC] = 8'h00;
mem[16'h3FBD] = 8'h00;
mem[16'h3FBE] = 8'h00;
mem[16'h3FBF] = 8'h00;
mem[16'h3FC0] = 8'h00;
mem[16'h3FC1] = 8'h00;
mem[16'h3FC2] = 8'h00;
mem[16'h3FC3] = 8'h00;
mem[16'h3FC4] = 8'h00;
mem[16'h3FC5] = 8'h00;
mem[16'h3FC6] = 8'h00;
mem[16'h3FC7] = 8'h00;
mem[16'h3FC8] = 8'h00;
mem[16'h3FC9] = 8'h00;
mem[16'h3FCA] = 8'h00;
mem[16'h3FCB] = 8'h00;
mem[16'h3FCC] = 8'h00;
mem[16'h3FCD] = 8'h00;
mem[16'h3FCE] = 8'h00;
mem[16'h3FCF] = 8'h2A;
mem[16'h3FD0] = 8'h00;
mem[16'h3FD1] = 8'h00;
mem[16'h3FD2] = 8'h00;
mem[16'h3FD3] = 8'h00;
mem[16'h3FD4] = 8'h00;
mem[16'h3FD5] = 8'h00;
mem[16'h3FD6] = 8'h00;
mem[16'h3FD7] = 8'h00;
mem[16'h3FD8] = 8'h00;
mem[16'h3FD9] = 8'h00;
mem[16'h3FDA] = 8'h00;
mem[16'h3FDB] = 8'h00;
mem[16'h3FDC] = 8'h00;
mem[16'h3FDD] = 8'h00;
mem[16'h3FDE] = 8'h00;
mem[16'h3FDF] = 8'h00;
mem[16'h3FE0] = 8'h00;
mem[16'h3FE1] = 8'h00;
mem[16'h3FE2] = 8'h00;
mem[16'h3FE3] = 8'h00;
mem[16'h3FE4] = 8'h00;
mem[16'h3FE5] = 8'h00;
mem[16'h3FE6] = 8'h00;
mem[16'h3FE7] = 8'h00;
mem[16'h3FE8] = 8'h00;
mem[16'h3FE9] = 8'h00;
mem[16'h3FEA] = 8'h00;
mem[16'h3FEB] = 8'h00;
mem[16'h3FEC] = 8'h00;
mem[16'h3FED] = 8'h00;
mem[16'h3FEE] = 8'h00;
mem[16'h3FEF] = 8'h00;
mem[16'h3FF0] = 8'h00;
mem[16'h3FF1] = 8'h00;
mem[16'h3FF2] = 8'h00;
mem[16'h3FF3] = 8'h00;
mem[16'h3FF4] = 8'h00;
mem[16'h3FF5] = 8'h00;
mem[16'h3FF6] = 8'h00;
mem[16'h3FF7] = 8'h00;
mem[16'h3FF8] = 8'h00;
mem[16'h3FF9] = 8'h00;
mem[16'h3FFA] = 8'h00;
mem[16'h3FFB] = 8'h00;
mem[16'h3FFC] = 8'h00;
mem[16'h3FFD] = 8'h00;
mem[16'h3FFE] = 8'h00;
mem[16'h3FFF] = 8'h00;
mem[16'h4000] = 8'h20;
mem[16'h4001] = 8'h83;
mem[16'h4002] = 8'h8B;
mem[16'h4003] = 8'h20;
mem[16'h4004] = 8'h00;
mem[16'h4005] = 8'h03;
mem[16'h4006] = 8'h20;
mem[16'h4007] = 8'h49;
mem[16'h4008] = 8'h71;
mem[16'h4009] = 8'h20;
mem[16'h400A] = 8'hCA;
mem[16'h400B] = 8'h5F;
mem[16'h400C] = 8'h20;
mem[16'h400D] = 8'h76;
mem[16'h400E] = 8'h41;
mem[16'h400F] = 8'h20;
mem[16'h4010] = 8'h42;
mem[16'h4011] = 8'h65;
mem[16'h4012] = 8'h20;
mem[16'h4013] = 8'h2F;
mem[16'h4014] = 8'h65;
mem[16'h4015] = 8'h6C;
mem[16'h4016] = 8'h5E;
mem[16'h4017] = 8'h00;
mem[16'h4018] = 8'h20;
mem[16'h4019] = 8'h96;
mem[16'h401A] = 8'h5D;
mem[16'h401B] = 8'h20;
mem[16'h401C] = 8'hA3;
mem[16'h401D] = 8'h55;
mem[16'h401E] = 8'h20;
mem[16'h401F] = 8'h25;
mem[16'h4020] = 8'h55;
mem[16'h4021] = 8'h20;
mem[16'h4022] = 8'h55;
mem[16'h4023] = 8'h90;
mem[16'h4024] = 8'h20;
mem[16'h4025] = 8'hCF;
mem[16'h4026] = 8'h44;
mem[16'h4027] = 8'h20;
mem[16'h4028] = 8'h2C;
mem[16'h4029] = 8'h53;
mem[16'h402A] = 8'h20;
mem[16'h402B] = 8'h9D;
mem[16'h402C] = 8'h51;
mem[16'h402D] = 8'h20;
mem[16'h402E] = 8'h97;
mem[16'h402F] = 8'h4F;
mem[16'h4030] = 8'h20;
mem[16'h4031] = 8'h05;
mem[16'h4032] = 8'h5E;
mem[16'h4033] = 8'h20;
mem[16'h4034] = 8'h64;
mem[16'h4035] = 8'h5E;
mem[16'h4036] = 8'h20;
mem[16'h4037] = 8'h36;
mem[16'h4038] = 8'h7B;
mem[16'h4039] = 8'h20;
mem[16'h403A] = 8'hFF;
mem[16'h403B] = 8'h44;
mem[16'h403C] = 8'h20;
mem[16'h403D] = 8'h62;
mem[16'h403E] = 8'h67;
mem[16'h403F] = 8'h20;
mem[16'h4040] = 8'h97;
mem[16'h4041] = 8'h90;
mem[16'h4042] = 8'h20;
mem[16'h4043] = 8'hB4;
mem[16'h4044] = 8'h4D;
mem[16'h4045] = 8'hA9;
mem[16'h4046] = 8'h17;
mem[16'h4047] = 8'h85;
mem[16'h4048] = 8'h25;
mem[16'h4049] = 8'hA9;
mem[16'h404A] = 8'h25;
mem[16'h404B] = 8'h85;
mem[16'h404C] = 8'h24;
mem[16'h404D] = 8'hAD;
mem[16'h404E] = 8'h50;
mem[16'h404F] = 8'h7F;
mem[16'h4050] = 8'h20;
mem[16'h4051] = 8'hED;
mem[16'h4052] = 8'hFD;
mem[16'h4053] = 8'h20;
mem[16'h4054] = 8'hC8;
mem[16'h4055] = 8'h6F;
mem[16'h4056] = 8'h20;
mem[16'h4057] = 8'hFC;
mem[16'h4058] = 8'h86;
mem[16'h4059] = 8'h20;
mem[16'h405A] = 8'h62;
mem[16'h405B] = 8'h5C;
mem[16'h405C] = 8'h20;
mem[16'h405D] = 8'hF7;
mem[16'h405E] = 8'h4F;
mem[16'h405F] = 8'h20;
mem[16'h4060] = 8'h28;
mem[16'h4061] = 8'h5C;
mem[16'h4062] = 8'h20;
mem[16'h4063] = 8'h43;
mem[16'h4064] = 8'h57;
mem[16'h4065] = 8'h20;
mem[16'h4066] = 8'h87;
mem[16'h4067] = 8'h58;
mem[16'h4068] = 8'h20;
mem[16'h4069] = 8'hFF;
mem[16'h406A] = 8'h55;
mem[16'h406B] = 8'h20;
mem[16'h406C] = 8'h63;
mem[16'h406D] = 8'h85;
mem[16'h406E] = 8'hA5;
mem[16'h406F] = 8'h73;
mem[16'h4070] = 8'hC9;
mem[16'h4071] = 8'h06;
mem[16'h4072] = 8'hD0;
mem[16'h4073] = 8'h06;
mem[16'h4074] = 8'h20;
mem[16'h4075] = 8'h62;
mem[16'h4076] = 8'h5C;
mem[16'h4077] = 8'h20;
mem[16'h4078] = 8'h43;
mem[16'h4079] = 8'h57;
mem[16'h407A] = 8'hAD;
mem[16'h407B] = 8'hB9;
mem[16'h407C] = 8'h4A;
mem[16'h407D] = 8'hC9;
mem[16'h407E] = 8'h02;
mem[16'h407F] = 8'h90;
mem[16'h4080] = 8'h03;
mem[16'h4081] = 8'h20;
mem[16'h4082] = 8'h28;
mem[16'h4083] = 8'h5C;
mem[16'h4084] = 8'hAD;
mem[16'h4085] = 8'hBA;
mem[16'h4086] = 8'h4A;
mem[16'h4087] = 8'hC9;
mem[16'h4088] = 8'h02;
mem[16'h4089] = 8'h90;
mem[16'h408A] = 8'h03;
mem[16'h408B] = 8'h20;
mem[16'h408C] = 8'h43;
mem[16'h408D] = 8'h57;
mem[16'h408E] = 8'h20;
mem[16'h408F] = 8'h18;
mem[16'h4090] = 8'h52;
mem[16'h4091] = 8'h20;
mem[16'h4092] = 8'hB4;
mem[16'h4093] = 8'h85;
mem[16'h4094] = 8'h20;
mem[16'h4095] = 8'hFB;
mem[16'h4096] = 8'h85;
mem[16'h4097] = 8'h20;
mem[16'h4098] = 8'hB0;
mem[16'h4099] = 8'h5A;
mem[16'h409A] = 8'h20;
mem[16'h409B] = 8'hE7;
mem[16'h409C] = 8'h59;
mem[16'h409D] = 8'h20;
mem[16'h409E] = 8'hDA;
mem[16'h409F] = 8'h77;
mem[16'h40A0] = 8'hAD;
mem[16'h40A1] = 8'hBA;
mem[16'h40A2] = 8'h4A;
mem[16'h40A3] = 8'hC9;
mem[16'h40A4] = 8'h03;
mem[16'h40A5] = 8'h90;
mem[16'h40A6] = 8'h03;
mem[16'h40A7] = 8'h20;
mem[16'h40A8] = 8'h43;
mem[16'h40A9] = 8'h57;
mem[16'h40AA] = 8'hAD;
mem[16'h40AB] = 8'hB8;
mem[16'h40AC] = 8'h4A;
mem[16'h40AD] = 8'hC9;
mem[16'h40AE] = 8'h02;
mem[16'h40AF] = 8'h90;
mem[16'h40B0] = 8'h03;
mem[16'h40B1] = 8'h20;
mem[16'h40B2] = 8'hFF;
mem[16'h40B3] = 8'h55;
mem[16'h40B4] = 8'h20;
mem[16'h40B5] = 8'hBD;
mem[16'h40B6] = 8'h4A;
mem[16'h40B7] = 8'h20;
mem[16'h40B8] = 8'h36;
mem[16'h40B9] = 8'h73;
mem[16'h40BA] = 8'h20;
mem[16'h40BB] = 8'h8A;
mem[16'h40BC] = 8'h53;
mem[16'h40BD] = 8'h20;
mem[16'h40BE] = 8'h35;
mem[16'h40BF] = 8'h45;
mem[16'h40C0] = 8'h20;
mem[16'h40C1] = 8'h48;
mem[16'h40C2] = 8'h47;
mem[16'h40C3] = 8'h20;
mem[16'h40C4] = 8'hD3;
mem[16'h40C5] = 8'h41;
mem[16'h40C6] = 8'h20;
mem[16'h40C7] = 8'hDD;
mem[16'h40C8] = 8'h42;
mem[16'h40C9] = 8'h20;
mem[16'h40CA] = 8'h09;
mem[16'h40CB] = 8'h6B;
mem[16'h40CC] = 8'h20;
mem[16'h40CD] = 8'h55;
mem[16'h40CE] = 8'h6A;
mem[16'h40CF] = 8'hAD;
mem[16'h40D0] = 8'hB9;
mem[16'h40D1] = 8'h4A;
mem[16'h40D2] = 8'hC9;
mem[16'h40D3] = 8'h03;
mem[16'h40D4] = 8'h90;
mem[16'h40D5] = 8'h03;
mem[16'h40D6] = 8'h20;
mem[16'h40D7] = 8'h28;
mem[16'h40D8] = 8'h5C;
mem[16'h40D9] = 8'hAD;
mem[16'h40DA] = 8'hB5;
mem[16'h40DB] = 8'h4A;
mem[16'h40DC] = 8'hC9;
mem[16'h40DD] = 8'h02;
mem[16'h40DE] = 8'h90;
mem[16'h40DF] = 8'h1C;
mem[16'h40E0] = 8'h20;
mem[16'h40E1] = 8'hF7;
mem[16'h40E2] = 8'h4F;
mem[16'h40E3] = 8'hA9;
mem[16'h40E4] = 8'h01;
mem[16'h40E5] = 8'h85;
mem[16'h40E6] = 8'h8B;
mem[16'h40E7] = 8'h20;
mem[16'h40E8] = 8'h09;
mem[16'h40E9] = 8'h6B;
mem[16'h40EA] = 8'h20;
mem[16'h40EB] = 8'h55;
mem[16'h40EC] = 8'h6A;
mem[16'h40ED] = 8'hA9;
mem[16'h40EE] = 8'h00;
mem[16'h40EF] = 8'h85;
mem[16'h40F0] = 8'h8B;
mem[16'h40F1] = 8'hAD;
mem[16'h40F2] = 8'h63;
mem[16'h40F3] = 8'h79;
mem[16'h40F4] = 8'hCD;
mem[16'h40F5] = 8'h13;
mem[16'h40F6] = 8'h51;
mem[16'h40F7] = 8'hD0;
mem[16'h40F8] = 8'h03;
mem[16'h40F9] = 8'h20;
mem[16'h40FA] = 8'hDA;
mem[16'h40FB] = 8'h77;
mem[16'h40FC] = 8'hAD;
mem[16'h40FD] = 8'hB6;
mem[16'h40FE] = 8'h4A;
mem[16'h40FF] = 8'hC9;
mem[16'h4100] = 8'h02;
mem[16'h4101] = 8'h90;
mem[16'h4102] = 8'h0E;
mem[16'h4103] = 8'h20;
mem[16'h4104] = 8'hE7;
mem[16'h4105] = 8'h59;
mem[16'h4106] = 8'hAD;
mem[16'h4107] = 8'h63;
mem[16'h4108] = 8'h79;
mem[16'h4109] = 8'hCD;
mem[16'h410A] = 8'h26;
mem[16'h410B] = 8'h5F;
mem[16'h410C] = 8'hD0;
mem[16'h410D] = 8'h03;
mem[16'h410E] = 8'h20;
mem[16'h410F] = 8'hDA;
mem[16'h4110] = 8'h77;
mem[16'h4111] = 8'hAD;
mem[16'h4112] = 8'hB4;
mem[16'h4113] = 8'h4A;
mem[16'h4114] = 8'hC9;
mem[16'h4115] = 8'h02;
mem[16'h4116] = 8'h90;
mem[16'h4117] = 8'h17;
mem[16'h4118] = 8'hA5;
mem[16'h4119] = 8'h73;
mem[16'h411A] = 8'h29;
mem[16'h411B] = 8'h01;
mem[16'h411C] = 8'hD0;
mem[16'h411D] = 8'h11;
mem[16'h411E] = 8'h20;
mem[16'h411F] = 8'h8A;
mem[16'h4120] = 8'h53;
mem[16'h4121] = 8'h20;
mem[16'h4122] = 8'h36;
mem[16'h4123] = 8'h73;
mem[16'h4124] = 8'hAD;
mem[16'h4125] = 8'h63;
mem[16'h4126] = 8'h79;
mem[16'h4127] = 8'hCD;
mem[16'h4128] = 8'h03;
mem[16'h4129] = 8'h54;
mem[16'h412A] = 8'hD0;
mem[16'h412B] = 8'h03;
mem[16'h412C] = 8'h20;
mem[16'h412D] = 8'hDA;
mem[16'h412E] = 8'h77;
mem[16'h412F] = 8'hAD;
mem[16'h4130] = 8'hB7;
mem[16'h4131] = 8'h4A;
mem[16'h4132] = 8'hC9;
mem[16'h4133] = 8'h02;
mem[16'h4134] = 8'hD0;
mem[16'h4135] = 8'h11;
mem[16'h4136] = 8'h20;
mem[16'h4137] = 8'hB0;
mem[16'h4138] = 8'h5A;
mem[16'h4139] = 8'hAD;
mem[16'h413A] = 8'h63;
mem[16'h413B] = 8'h79;
mem[16'h413C] = 8'hCD;
mem[16'h413D] = 8'h1E;
mem[16'h413E] = 8'h5F;
mem[16'h413F] = 8'hD0;
mem[16'h4140] = 8'h1A;
mem[16'h4141] = 8'h20;
mem[16'h4142] = 8'hDA;
mem[16'h4143] = 8'h77;
mem[16'h4144] = 8'h4C;
mem[16'h4145] = 8'h5B;
mem[16'h4146] = 8'h41;
mem[16'h4147] = 8'hA5;
mem[16'h4148] = 8'h73;
mem[16'h4149] = 8'h29;
mem[16'h414A] = 8'h01;
mem[16'h414B] = 8'hD0;
mem[16'h414C] = 8'h0E;
mem[16'h414D] = 8'h20;
mem[16'h414E] = 8'hB0;
mem[16'h414F] = 8'h5A;
mem[16'h4150] = 8'hAD;
mem[16'h4151] = 8'h63;
mem[16'h4152] = 8'h79;
mem[16'h4153] = 8'hCD;
mem[16'h4154] = 8'h1E;
mem[16'h4155] = 8'h5F;
mem[16'h4156] = 8'hD0;
mem[16'h4157] = 8'h03;
mem[16'h4158] = 8'h20;
mem[16'h4159] = 8'hDA;
mem[16'h415A] = 8'h77;
mem[16'h415B] = 8'hA5;
mem[16'h415C] = 8'h73;
mem[16'h415D] = 8'h29;
mem[16'h415E] = 8'h01;
mem[16'h415F] = 8'hF0;
mem[16'h4160] = 8'h03;
mem[16'h4161] = 8'h20;
mem[16'h4162] = 8'hDA;
mem[16'h4163] = 8'h77;
mem[16'h4164] = 8'h20;
mem[16'h4165] = 8'hD4;
mem[16'h4166] = 8'h90;
mem[16'h4167] = 8'h20;
mem[16'h4168] = 8'hD0;
mem[16'h4169] = 8'h7F;
mem[16'h416A] = 8'h20;
mem[16'h416B] = 8'h01;
mem[16'h416C] = 8'h7F;
mem[16'h416D] = 8'h20;
mem[16'h416E] = 8'hF1;
mem[16'h416F] = 8'h6F;
mem[16'h4170] = 8'h20;
mem[16'h4171] = 8'hDC;
mem[16'h4172] = 8'h6F;
mem[16'h4173] = 8'h4C;
mem[16'h4174] = 8'h56;
mem[16'h4175] = 8'h40;
mem[16'h4176] = 8'hA9;
mem[16'h4177] = 8'h00;
mem[16'h4178] = 8'h8D;
mem[16'h4179] = 8'hD2;
mem[16'h417A] = 8'h67;
mem[16'h417B] = 8'h8D;
mem[16'h417C] = 8'hD3;
mem[16'h417D] = 8'h67;
mem[16'h417E] = 8'h8D;
mem[16'h417F] = 8'hD4;
mem[16'h4180] = 8'h67;
mem[16'h4181] = 8'h8D;
mem[16'h4182] = 8'hCF;
mem[16'h4183] = 8'h67;
mem[16'h4184] = 8'h8D;
mem[16'h4185] = 8'hD0;
mem[16'h4186] = 8'h67;
mem[16'h4187] = 8'h8D;
mem[16'h4188] = 8'hD1;
mem[16'h4189] = 8'h67;
mem[16'h418A] = 8'hA9;
mem[16'h418B] = 8'h01;
mem[16'h418C] = 8'h8D;
mem[16'h418D] = 8'hCD;
mem[16'h418E] = 8'h6A;
mem[16'h418F] = 8'h8D;
mem[16'h4190] = 8'h88;
mem[16'h4191] = 8'h6B;
mem[16'h4192] = 8'hA9;
mem[16'h4193] = 8'h5E;
mem[16'h4194] = 8'h8D;
mem[16'h4195] = 8'hC9;
mem[16'h4196] = 8'h77;
mem[16'h4197] = 8'h8D;
mem[16'h4198] = 8'hCB;
mem[16'h4199] = 8'h77;
mem[16'h419A] = 8'hA9;
mem[16'h419B] = 8'h06;
mem[16'h419C] = 8'h8D;
mem[16'h419D] = 8'hE0;
mem[16'h419E] = 8'h91;
mem[16'h419F] = 8'hAD;
mem[16'h41A0] = 8'h14;
mem[16'h41A1] = 8'h87;
mem[16'h41A2] = 8'h29;
mem[16'h41A3] = 8'h3F;
mem[16'h41A4] = 8'h8D;
mem[16'h41A5] = 8'hD8;
mem[16'h41A6] = 8'h91;
mem[16'h41A7] = 8'hA9;
mem[16'h41A8] = 8'hC8;
mem[16'h41A9] = 8'h8D;
mem[16'h41AA] = 8'hD9;
mem[16'h41AB] = 8'h91;
mem[16'h41AC] = 8'hA9;
mem[16'h41AD] = 8'h01;
mem[16'h41AE] = 8'h8D;
mem[16'h41AF] = 8'hCE;
mem[16'h41B0] = 8'h44;
mem[16'h41B1] = 8'hA9;
mem[16'h41B2] = 8'h05;
mem[16'h41B3] = 8'h8D;
mem[16'h41B4] = 8'hE6;
mem[16'h41B5] = 8'h48;
mem[16'h41B6] = 8'hA9;
mem[16'h41B7] = 8'h55;
mem[16'h41B8] = 8'h85;
mem[16'h41B9] = 8'h5E;
mem[16'h41BA] = 8'hA9;
mem[16'h41BB] = 8'h49;
mem[16'h41BC] = 8'h85;
mem[16'h41BD] = 8'h5F;
mem[16'h41BE] = 8'hA9;
mem[16'h41BF] = 8'h00;
mem[16'h41C0] = 8'h8D;
mem[16'h41C1] = 8'hA8;
mem[16'h41C2] = 8'h44;
mem[16'h41C3] = 8'h8D;
mem[16'h41C4] = 8'h5E;
mem[16'h41C5] = 8'h42;
mem[16'h41C6] = 8'h8D;
mem[16'h41C7] = 8'h5F;
mem[16'h41C8] = 8'h42;
mem[16'h41C9] = 8'h8D;
mem[16'h41CA] = 8'h60;
mem[16'h41CB] = 8'h42;
mem[16'h41CC] = 8'h8D;
mem[16'h41CD] = 8'h61;
mem[16'h41CE] = 8'h42;
mem[16'h41CF] = 8'h8D;
mem[16'h41D0] = 8'h62;
mem[16'h41D1] = 8'h42;
mem[16'h41D2] = 8'h60;
mem[16'h41D3] = 8'hCE;
mem[16'h41D4] = 8'h57;
mem[16'h41D5] = 8'h42;
mem[16'h41D6] = 8'hF0;
mem[16'h41D7] = 8'h2C;
mem[16'h41D8] = 8'hAD;
mem[16'h41D9] = 8'h57;
mem[16'h41DA] = 8'h42;
mem[16'h41DB] = 8'hC9;
mem[16'h41DC] = 8'hFC;
mem[16'h41DD] = 8'hF0;
mem[16'h41DE] = 8'h48;
mem[16'h41DF] = 8'hC9;
mem[16'h41E0] = 8'hF9;
mem[16'h41E1] = 8'hF0;
mem[16'h41E2] = 8'h5C;
mem[16'h41E3] = 8'hC9;
mem[16'h41E4] = 8'hB4;
mem[16'h41E5] = 8'hD0;
mem[16'h41E6] = 8'h13;
mem[16'h41E7] = 8'hAE;
mem[16'h41E8] = 8'h58;
mem[16'h41E9] = 8'h42;
mem[16'h41EA] = 8'hBD;
mem[16'h41EB] = 8'h5E;
mem[16'h41EC] = 8'h42;
mem[16'h41ED] = 8'hC9;
mem[16'h41EE] = 8'h03;
mem[16'h41EF] = 8'hD0;
mem[16'h41F0] = 8'h12;
mem[16'h41F1] = 8'hA9;
mem[16'h41F2] = 8'h00;
mem[16'h41F3] = 8'h9D;
mem[16'h41F4] = 8'h5E;
mem[16'h41F5] = 8'h42;
mem[16'h41F6] = 8'h20;
mem[16'h41F7] = 8'h63;
mem[16'h41F8] = 8'h42;
mem[16'h41F9] = 8'h60;
mem[16'h41FA] = 8'hC9;
mem[16'h41FB] = 8'h32;
mem[16'h41FC] = 8'hD0;
mem[16'h41FD] = 8'h05;
mem[16'h41FE] = 8'hA9;
mem[16'h41FF] = 8'h01;
mem[16'h4200] = 8'h8D;
mem[16'h4201] = 8'h57;
mem[16'h4202] = 8'h42;
mem[16'h4203] = 8'h60;
mem[16'h4204] = 8'hAE;
mem[16'h4205] = 8'h58;
mem[16'h4206] = 8'h42;
mem[16'h4207] = 8'hCA;
mem[16'h4208] = 8'h10;
mem[16'h4209] = 8'h02;
mem[16'h420A] = 8'hA2;
mem[16'h420B] = 8'h04;
mem[16'h420C] = 8'h8E;
mem[16'h420D] = 8'h58;
mem[16'h420E] = 8'h42;
mem[16'h420F] = 8'hBD;
mem[16'h4210] = 8'h5E;
mem[16'h4211] = 8'h42;
mem[16'h4212] = 8'hD0;
mem[16'h4213] = 8'hEF;
mem[16'h4214] = 8'hBD;
mem[16'h4215] = 8'h59;
mem[16'h4216] = 8'h42;
mem[16'h4217] = 8'h8D;
mem[16'h4218] = 8'h8F;
mem[16'h4219] = 8'h42;
mem[16'h421A] = 8'hA9;
mem[16'h421B] = 8'h03;
mem[16'h421C] = 8'h9D;
mem[16'h421D] = 8'h5E;
mem[16'h421E] = 8'h42;
mem[16'h421F] = 8'hA9;
mem[16'h4220] = 8'hA7;
mem[16'h4221] = 8'hA0;
mem[16'h4222] = 8'h42;
mem[16'h4223] = 8'h20;
mem[16'h4224] = 8'h91;
mem[16'h4225] = 8'h42;
mem[16'h4226] = 8'h60;
mem[16'h4227] = 8'hAE;
mem[16'h4228] = 8'h58;
mem[16'h4229] = 8'h42;
mem[16'h422A] = 8'hBD;
mem[16'h422B] = 8'h5E;
mem[16'h422C] = 8'h42;
mem[16'h422D] = 8'hC9;
mem[16'h422E] = 8'h03;
mem[16'h422F] = 8'hD0;
mem[16'h4230] = 8'hD2;
mem[16'h4231] = 8'hBD;
mem[16'h4232] = 8'h59;
mem[16'h4233] = 8'h42;
mem[16'h4234] = 8'h8D;
mem[16'h4235] = 8'h8F;
mem[16'h4236] = 8'h42;
mem[16'h4237] = 8'hA9;
mem[16'h4238] = 8'hB9;
mem[16'h4239] = 8'hA0;
mem[16'h423A] = 8'h42;
mem[16'h423B] = 8'h20;
mem[16'h423C] = 8'h91;
mem[16'h423D] = 8'h42;
mem[16'h423E] = 8'h60;
mem[16'h423F] = 8'hAE;
mem[16'h4240] = 8'h58;
mem[16'h4241] = 8'h42;
mem[16'h4242] = 8'hBD;
mem[16'h4243] = 8'h5E;
mem[16'h4244] = 8'h42;
mem[16'h4245] = 8'hC9;
mem[16'h4246] = 8'h03;
mem[16'h4247] = 8'hD0;
mem[16'h4248] = 8'hBA;
mem[16'h4249] = 8'hBD;
mem[16'h424A] = 8'h59;
mem[16'h424B] = 8'h42;
mem[16'h424C] = 8'h8D;
mem[16'h424D] = 8'h8F;
mem[16'h424E] = 8'h42;
mem[16'h424F] = 8'hA9;
mem[16'h4250] = 8'hCB;
mem[16'h4251] = 8'hA0;
mem[16'h4252] = 8'h42;
mem[16'h4253] = 8'h20;
mem[16'h4254] = 8'h91;
mem[16'h4255] = 8'h42;
mem[16'h4256] = 8'h60;
mem[16'h4257] = 8'hB4;
mem[16'h4258] = 8'h02;
mem[16'h4259] = 8'h46;
mem[16'h425A] = 8'hCC;
mem[16'h425B] = 8'h16;
mem[16'h425C] = 8'hA2;
mem[16'h425D] = 8'h70;
mem[16'h425E] = 8'h00;
mem[16'h425F] = 8'h00;
mem[16'h4260] = 8'h00;
mem[16'h4261] = 8'h00;
mem[16'h4262] = 8'h00;
mem[16'h4263] = 8'hA9;
mem[16'h4264] = 8'h7D;
mem[16'h4265] = 8'hA0;
mem[16'h4266] = 8'h42;
mem[16'h4267] = 8'h20;
mem[16'h4268] = 8'h2B;
mem[16'h4269] = 8'h8C;
mem[16'h426A] = 8'hA9;
mem[16'h426B] = 8'h12;
mem[16'h426C] = 8'h8D;
mem[16'h426D] = 8'h24;
mem[16'h426E] = 8'h8C;
mem[16'h426F] = 8'hAD;
mem[16'h4270] = 8'h8F;
mem[16'h4271] = 8'h42;
mem[16'h4272] = 8'h85;
mem[16'h4273] = 8'h57;
mem[16'h4274] = 8'hAD;
mem[16'h4275] = 8'h90;
mem[16'h4276] = 8'h42;
mem[16'h4277] = 8'h85;
mem[16'h4278] = 8'h56;
mem[16'h4279] = 8'h20;
mem[16'h427A] = 8'hA8;
mem[16'h427B] = 8'h8B;
mem[16'h427C] = 8'h60;
mem[16'h427D] = 8'h55;
mem[16'h427E] = 8'h2A;
mem[16'h427F] = 8'h5F;
mem[16'h4280] = 8'h3E;
mem[16'h4281] = 8'h57;
mem[16'h4282] = 8'h3F;
mem[16'h4283] = 8'h7F;
mem[16'h4284] = 8'h2B;
mem[16'h4285] = 8'h57;
mem[16'h4286] = 8'h2A;
mem[16'h4287] = 8'h7F;
mem[16'h4288] = 8'h3F;
mem[16'h4289] = 8'h7F;
mem[16'h428A] = 8'h3F;
mem[16'h428B] = 8'h7F;
mem[16'h428C] = 8'h2A;
mem[16'h428D] = 8'h55;
mem[16'h428E] = 8'h2A;
mem[16'h428F] = 8'h85;
mem[16'h4290] = 8'h0A;
mem[16'h4291] = 8'h20;
mem[16'h4292] = 8'h2B;
mem[16'h4293] = 8'h8C;
mem[16'h4294] = 8'hA9;
mem[16'h4295] = 8'h12;
mem[16'h4296] = 8'h8D;
mem[16'h4297] = 8'h24;
mem[16'h4298] = 8'h8C;
mem[16'h4299] = 8'hAD;
mem[16'h429A] = 8'h8F;
mem[16'h429B] = 8'h42;
mem[16'h429C] = 8'h85;
mem[16'h429D] = 8'h57;
mem[16'h429E] = 8'hAD;
mem[16'h429F] = 8'h90;
mem[16'h42A0] = 8'h42;
mem[16'h42A1] = 8'h85;
mem[16'h42A2] = 8'h56;
mem[16'h42A3] = 8'h20;
mem[16'h42A4] = 8'hA8;
mem[16'h42A5] = 8'h8B;
mem[16'h42A6] = 8'h60;
mem[16'h42A7] = 8'h55;
mem[16'h42A8] = 8'h2A;
mem[16'h42A9] = 8'h57;
mem[16'h42AA] = 8'h2E;
mem[16'h42AB] = 8'h55;
mem[16'h42AC] = 8'h3B;
mem[16'h42AD] = 8'h75;
mem[16'h42AE] = 8'h2A;
mem[16'h42AF] = 8'h57;
mem[16'h42B0] = 8'h2A;
mem[16'h42B1] = 8'h55;
mem[16'h42B2] = 8'h2E;
mem[16'h42B3] = 8'h5D;
mem[16'h42B4] = 8'h2A;
mem[16'h42B5] = 8'h75;
mem[16'h42B6] = 8'h2A;
mem[16'h42B7] = 8'h55;
mem[16'h42B8] = 8'h2A;
mem[16'h42B9] = 8'h00;
mem[16'h42BA] = 8'h00;
mem[16'h42BB] = 8'h08;
mem[16'h42BC] = 8'h00;
mem[16'h42BD] = 8'h00;
mem[16'h42BE] = 8'h00;
mem[16'h42BF] = 8'h02;
mem[16'h42C0] = 8'h00;
mem[16'h42C1] = 8'h00;
mem[16'h42C2] = 8'h00;
mem[16'h42C3] = 8'h28;
mem[16'h42C4] = 8'h10;
mem[16'h42C5] = 8'h00;
mem[16'h42C6] = 8'h01;
mem[16'h42C7] = 8'h02;
mem[16'h42C8] = 8'h00;
mem[16'h42C9] = 8'h00;
mem[16'h42CA] = 8'h00;
mem[16'h42CB] = 8'h00;
mem[16'h42CC] = 8'h00;
mem[16'h42CD] = 8'h00;
mem[16'h42CE] = 8'h10;
mem[16'h42CF] = 8'h02;
mem[16'h42D0] = 8'h04;
mem[16'h42D1] = 8'h08;
mem[16'h42D2] = 8'h01;
mem[16'h42D3] = 8'h00;
mem[16'h42D4] = 8'h00;
mem[16'h42D5] = 8'h02;
mem[16'h42D6] = 8'h01;
mem[16'h42D7] = 8'h22;
mem[16'h42D8] = 8'h14;
mem[16'h42D9] = 8'h08;
mem[16'h42DA] = 8'h00;
mem[16'h42DB] = 8'h00;
mem[16'h42DC] = 8'h00;
mem[16'h42DD] = 8'hCE;
mem[16'h42DE] = 8'h22;
mem[16'h42DF] = 8'h43;
mem[16'h42E0] = 8'hF0;
mem[16'h42E1] = 8'h1F;
mem[16'h42E2] = 8'hAD;
mem[16'h42E3] = 8'h22;
mem[16'h42E4] = 8'h43;
mem[16'h42E5] = 8'hC9;
mem[16'h42E6] = 8'h96;
mem[16'h42E7] = 8'hD0;
mem[16'h42E8] = 8'h17;
mem[16'h42E9] = 8'hA9;
mem[16'h42EA] = 8'h50;
mem[16'h42EB] = 8'h8D;
mem[16'h42EC] = 8'h22;
mem[16'h42ED] = 8'h43;
mem[16'h42EE] = 8'hAE;
mem[16'h42EF] = 8'h23;
mem[16'h42F0] = 8'h43;
mem[16'h42F1] = 8'hBD;
mem[16'h42F2] = 8'h5E;
mem[16'h42F3] = 8'h42;
mem[16'h42F4] = 8'hC9;
mem[16'h42F5] = 8'h02;
mem[16'h42F6] = 8'hD0;
mem[16'h42F7] = 8'h08;
mem[16'h42F8] = 8'hA9;
mem[16'h42F9] = 8'h00;
mem[16'h42FA] = 8'h9D;
mem[16'h42FB] = 8'h5E;
mem[16'h42FC] = 8'h42;
mem[16'h42FD] = 8'h20;
mem[16'h42FE] = 8'h29;
mem[16'h42FF] = 8'h43;
mem[16'h4300] = 8'h60;
mem[16'h4301] = 8'hAE;
mem[16'h4302] = 8'h23;
mem[16'h4303] = 8'h43;
mem[16'h4304] = 8'hE8;
mem[16'h4305] = 8'hE0;
mem[16'h4306] = 8'h05;
mem[16'h4307] = 8'h90;
mem[16'h4308] = 8'h02;
mem[16'h4309] = 8'hA2;
mem[16'h430A] = 8'h00;
mem[16'h430B] = 8'h8E;
mem[16'h430C] = 8'h23;
mem[16'h430D] = 8'h43;
mem[16'h430E] = 8'hBD;
mem[16'h430F] = 8'h5E;
mem[16'h4310] = 8'h42;
mem[16'h4311] = 8'hD0;
mem[16'h4312] = 8'hED;
mem[16'h4313] = 8'hBD;
mem[16'h4314] = 8'h24;
mem[16'h4315] = 8'h43;
mem[16'h4316] = 8'h8D;
mem[16'h4317] = 8'h57;
mem[16'h4318] = 8'h43;
mem[16'h4319] = 8'hA9;
mem[16'h431A] = 8'h02;
mem[16'h431B] = 8'h9D;
mem[16'h431C] = 8'h5E;
mem[16'h431D] = 8'h42;
mem[16'h431E] = 8'h20;
mem[16'h431F] = 8'h29;
mem[16'h4320] = 8'h43;
mem[16'h4321] = 8'h60;
mem[16'h4322] = 8'hC8;
mem[16'h4323] = 8'h01;
mem[16'h4324] = 8'h46;
mem[16'h4325] = 8'hCA;
mem[16'h4326] = 8'h14;
mem[16'h4327] = 8'hA0;
mem[16'h4328] = 8'h70;
mem[16'h4329] = 8'hA9;
mem[16'h432A] = 8'h43;
mem[16'h432B] = 8'hA0;
mem[16'h432C] = 8'h43;
mem[16'h432D] = 8'h20;
mem[16'h432E] = 8'h2B;
mem[16'h432F] = 8'h8C;
mem[16'h4330] = 8'hA9;
mem[16'h4331] = 8'h14;
mem[16'h4332] = 8'h8D;
mem[16'h4333] = 8'h24;
mem[16'h4334] = 8'h8C;
mem[16'h4335] = 8'hAD;
mem[16'h4336] = 8'h57;
mem[16'h4337] = 8'h43;
mem[16'h4338] = 8'h85;
mem[16'h4339] = 8'h57;
mem[16'h433A] = 8'hAD;
mem[16'h433B] = 8'h58;
mem[16'h433C] = 8'h43;
mem[16'h433D] = 8'h85;
mem[16'h433E] = 8'h56;
mem[16'h433F] = 8'h20;
mem[16'h4340] = 8'hA8;
mem[16'h4341] = 8'h8B;
mem[16'h4342] = 8'h60;
mem[16'h4343] = 8'h15;
mem[16'h4344] = 8'h2B;
mem[16'h4345] = 8'h35;
mem[16'h4346] = 8'h29;
mem[16'h4347] = 8'h15;
mem[16'h4348] = 8'h2B;
mem[16'h4349] = 8'h35;
mem[16'h434A] = 8'h29;
mem[16'h434B] = 8'h05;
mem[16'h434C] = 8'h2F;
mem[16'h434D] = 8'h0D;
mem[16'h434E] = 8'h27;
mem[16'h434F] = 8'h01;
mem[16'h4350] = 8'h3F;
mem[16'h4351] = 8'h61;
mem[16'h4352] = 8'h3C;
mem[16'h4353] = 8'h41;
mem[16'h4354] = 8'h3E;
mem[16'h4355] = 8'h59;
mem[16'h4356] = 8'h22;
mem[16'h4357] = 8'h09;
mem[16'h4358] = 8'h0A;
mem[16'h4359] = 8'hAD;
mem[16'h435A] = 8'hD0;
mem[16'h435B] = 8'h4D;
mem[16'h435C] = 8'hC9;
mem[16'h435D] = 8'h07;
mem[16'h435E] = 8'hF0;
mem[16'h435F] = 8'h01;
mem[16'h4360] = 8'h60;
mem[16'h4361] = 8'hAD;
mem[16'h4362] = 8'hCF;
mem[16'h4363] = 8'h4D;
mem[16'h4364] = 8'hA2;
mem[16'h4365] = 8'h02;
mem[16'h4366] = 8'h38;
mem[16'h4367] = 8'hE9;
mem[16'h4368] = 8'h15;
mem[16'h4369] = 8'h20;
mem[16'h436A] = 8'h62;
mem[16'h436B] = 8'h65;
mem[16'h436C] = 8'hC9;
mem[16'h436D] = 8'h04;
mem[16'h436E] = 8'h90;
mem[16'h436F] = 8'h3F;
mem[16'h4370] = 8'hA2;
mem[16'h4371] = 8'h00;
mem[16'h4372] = 8'hAD;
mem[16'h4373] = 8'hCF;
mem[16'h4374] = 8'h4D;
mem[16'h4375] = 8'h38;
mem[16'h4376] = 8'hE9;
mem[16'h4377] = 8'h46;
mem[16'h4378] = 8'h20;
mem[16'h4379] = 8'h62;
mem[16'h437A] = 8'h65;
mem[16'h437B] = 8'hC9;
mem[16'h437C] = 8'h04;
mem[16'h437D] = 8'h90;
mem[16'h437E] = 8'h30;
mem[16'h437F] = 8'hA2;
mem[16'h4380] = 8'h04;
mem[16'h4381] = 8'hAD;
mem[16'h4382] = 8'hCF;
mem[16'h4383] = 8'h4D;
mem[16'h4384] = 8'h38;
mem[16'h4385] = 8'hE9;
mem[16'h4386] = 8'h70;
mem[16'h4387] = 8'h20;
mem[16'h4388] = 8'h62;
mem[16'h4389] = 8'h65;
mem[16'h438A] = 8'hC9;
mem[16'h438B] = 8'h04;
mem[16'h438C] = 8'h90;
mem[16'h438D] = 8'h21;
mem[16'h438E] = 8'hA2;
mem[16'h438F] = 8'h03;
mem[16'h4390] = 8'hAD;
mem[16'h4391] = 8'hCF;
mem[16'h4392] = 8'h4D;
mem[16'h4393] = 8'h38;
mem[16'h4394] = 8'hE9;
mem[16'h4395] = 8'hA1;
mem[16'h4396] = 8'h20;
mem[16'h4397] = 8'h62;
mem[16'h4398] = 8'h65;
mem[16'h4399] = 8'hC9;
mem[16'h439A] = 8'h04;
mem[16'h439B] = 8'h90;
mem[16'h439C] = 8'h12;
mem[16'h439D] = 8'hA2;
mem[16'h439E] = 8'h01;
mem[16'h439F] = 8'hAD;
mem[16'h43A0] = 8'hCF;
mem[16'h43A1] = 8'h4D;
mem[16'h43A2] = 8'h38;
mem[16'h43A3] = 8'hE9;
mem[16'h43A4] = 8'hCB;
mem[16'h43A5] = 8'h20;
mem[16'h43A6] = 8'h62;
mem[16'h43A7] = 8'h65;
mem[16'h43A8] = 8'hC9;
mem[16'h43A9] = 8'h04;
mem[16'h43AA] = 8'h90;
mem[16'h43AB] = 8'h03;
mem[16'h43AC] = 8'h4C;
mem[16'h43AD] = 8'h8E;
mem[16'h43AE] = 8'h48;
mem[16'h43AF] = 8'hA9;
mem[16'h43B0] = 8'h00;
mem[16'h43B1] = 8'h8D;
mem[16'h43B2] = 8'h91;
mem[16'h43B3] = 8'h6F;
mem[16'h43B4] = 8'h8D;
mem[16'h43B5] = 8'hA9;
mem[16'h43B6] = 8'h44;
mem[16'h43B7] = 8'h86;
mem[16'h43B8] = 8'h70;
mem[16'h43B9] = 8'hBD;
mem[16'h43BA] = 8'h5E;
mem[16'h43BB] = 8'h42;
mem[16'h43BC] = 8'hC9;
mem[16'h43BD] = 8'h01;
mem[16'h43BE] = 8'hF0;
mem[16'h43BF] = 8'h0D;
mem[16'h43C0] = 8'hC9;
mem[16'h43C1] = 8'h03;
mem[16'h43C2] = 8'hD0;
mem[16'h43C3] = 8'h0C;
mem[16'h43C4] = 8'hAD;
mem[16'h43C5] = 8'h57;
mem[16'h43C6] = 8'h42;
mem[16'h43C7] = 8'hF0;
mem[16'h43C8] = 8'h07;
mem[16'h43C9] = 8'hC9;
mem[16'h43CA] = 8'hF9;
mem[16'h43CB] = 8'hB0;
mem[16'h43CC] = 8'h03;
mem[16'h43CD] = 8'h4C;
mem[16'h43CE] = 8'h8E;
mem[16'h43CF] = 8'h48;
mem[16'h43D0] = 8'hC9;
mem[16'h43D1] = 8'h02;
mem[16'h43D2] = 8'hD0;
mem[16'h43D3] = 8'h17;
mem[16'h43D4] = 8'hA9;
mem[16'h43D5] = 8'h02;
mem[16'h43D6] = 8'h20;
mem[16'h43D7] = 8'hAD;
mem[16'h43D8] = 8'h66;
mem[16'h43D9] = 8'hA6;
mem[16'h43DA] = 8'h70;
mem[16'h43DB] = 8'hBD;
mem[16'h43DC] = 8'hA3;
mem[16'h43DD] = 8'h44;
mem[16'h43DE] = 8'h18;
mem[16'h43DF] = 8'h69;
mem[16'h43E0] = 8'h12;
mem[16'h43E1] = 8'h09;
mem[16'h43E2] = 8'h01;
mem[16'h43E3] = 8'h8D;
mem[16'h43E4] = 8'h91;
mem[16'h43E5] = 8'h6F;
mem[16'h43E6] = 8'hEE;
mem[16'h43E7] = 8'hA9;
mem[16'h43E8] = 8'h44;
mem[16'h43E9] = 8'hA6;
mem[16'h43EA] = 8'h70;
mem[16'h43EB] = 8'hAD;
mem[16'h43EC] = 8'hB2;
mem[16'h43ED] = 8'h85;
mem[16'h43EE] = 8'hD0;
mem[16'h43EF] = 8'h06;
mem[16'h43F0] = 8'hAD;
mem[16'h43F1] = 8'hB1;
mem[16'h43F2] = 8'h85;
mem[16'h43F3] = 8'h8D;
mem[16'h43F4] = 8'hB0;
mem[16'h43F5] = 8'h85;
mem[16'h43F6] = 8'hAD;
mem[16'h43F7] = 8'hB3;
mem[16'h43F8] = 8'h85;
mem[16'h43F9] = 8'hF0;
mem[16'h43FA] = 8'h1F;
mem[16'h43FB] = 8'h86;
mem[16'h43FC] = 8'h70;
mem[16'h43FD] = 8'hA9;
mem[16'h43FE] = 8'h02;
mem[16'h43FF] = 8'h20;
mem[16'h4400] = 8'hAD;
mem[16'h4401] = 8'h66;
mem[16'h4402] = 8'h20;
mem[16'h4403] = 8'h0E;
mem[16'h4404] = 8'h73;
mem[16'h4405] = 8'hA9;
mem[16'h4406] = 8'h00;
mem[16'h4407] = 8'h8D;
mem[16'h4408] = 8'hB3;
mem[16'h4409] = 8'h85;
mem[16'h440A] = 8'hEE;
mem[16'h440B] = 8'hA9;
mem[16'h440C] = 8'h44;
mem[16'h440D] = 8'hA6;
mem[16'h440E] = 8'h70;
mem[16'h440F] = 8'hBD;
mem[16'h4410] = 8'hA3;
mem[16'h4411] = 8'h44;
mem[16'h4412] = 8'h18;
mem[16'h4413] = 8'h69;
mem[16'h4414] = 8'h12;
mem[16'h4415] = 8'h09;
mem[16'h4416] = 8'h01;
mem[16'h4417] = 8'h8D;
mem[16'h4418] = 8'h91;
mem[16'h4419] = 8'h6F;
mem[16'h441A] = 8'hAD;
mem[16'h441B] = 8'hA9;
mem[16'h441C] = 8'h44;
mem[16'h441D] = 8'hF0;
mem[16'h441E] = 8'h1C;
mem[16'h441F] = 8'hC9;
mem[16'h4420] = 8'h01;
mem[16'h4421] = 8'hF0;
mem[16'h4422] = 8'h07;
mem[16'h4423] = 8'hA9;
mem[16'h4424] = 8'hAD;
mem[16'h4425] = 8'hA0;
mem[16'h4426] = 8'h6F;
mem[16'h4427] = 8'h4C;
mem[16'h4428] = 8'h2E;
mem[16'h4429] = 8'h44;
mem[16'h442A] = 8'hA9;
mem[16'h442B] = 8'h92;
mem[16'h442C] = 8'hA0;
mem[16'h442D] = 8'h6F;
mem[16'h442E] = 8'h20;
mem[16'h442F] = 8'h86;
mem[16'h4430] = 8'h68;
mem[16'h4431] = 8'h85;
mem[16'h4432] = 8'h60;
mem[16'h4433] = 8'h84;
mem[16'h4434] = 8'h61;
mem[16'h4435] = 8'h20;
mem[16'h4436] = 8'hF8;
mem[16'h4437] = 8'h6E;
mem[16'h4438] = 8'h20;
mem[16'h4439] = 8'h23;
mem[16'h443A] = 8'h4C;
mem[16'h443B] = 8'hA6;
mem[16'h443C] = 8'h70;
mem[16'h443D] = 8'hA9;
mem[16'h443E] = 8'h01;
mem[16'h443F] = 8'hEE;
mem[16'h4440] = 8'hA8;
mem[16'h4441] = 8'h44;
mem[16'h4442] = 8'h9D;
mem[16'h4443] = 8'h5E;
mem[16'h4444] = 8'h42;
mem[16'h4445] = 8'h86;
mem[16'h4446] = 8'h70;
mem[16'h4447] = 8'h20;
mem[16'h4448] = 8'hD9;
mem[16'h4449] = 8'h4C;
mem[16'h444A] = 8'hA6;
mem[16'h444B] = 8'h70;
mem[16'h444C] = 8'hBD;
mem[16'h444D] = 8'hA3;
mem[16'h444E] = 8'h44;
mem[16'h444F] = 8'h8D;
mem[16'h4450] = 8'hCF;
mem[16'h4451] = 8'h4D;
mem[16'h4452] = 8'h20;
mem[16'h4453] = 8'hD9;
mem[16'h4454] = 8'h4C;
mem[16'h4455] = 8'hA9;
mem[16'h4456] = 8'h50;
mem[16'h4457] = 8'h20;
mem[16'h4458] = 8'h89;
mem[16'h4459] = 8'h66;
mem[16'h445A] = 8'h20;
mem[16'h445B] = 8'h43;
mem[16'h445C] = 8'h6E;
mem[16'h445D] = 8'hA9;
mem[16'h445E] = 8'h5A;
mem[16'h445F] = 8'h8D;
mem[16'h4460] = 8'h22;
mem[16'h4461] = 8'h4C;
mem[16'h4462] = 8'hA5;
mem[16'h4463] = 8'h74;
mem[16'h4464] = 8'h85;
mem[16'h4465] = 8'h72;
mem[16'h4466] = 8'hF8;
mem[16'h4467] = 8'hA5;
mem[16'h4468] = 8'h72;
mem[16'h4469] = 8'h38;
mem[16'h446A] = 8'hE9;
mem[16'h446B] = 8'h01;
mem[16'h446C] = 8'h85;
mem[16'h446D] = 8'h72;
mem[16'h446E] = 8'hF0;
mem[16'h446F] = 8'h0F;
mem[16'h4470] = 8'h30;
mem[16'h4471] = 8'h0D;
mem[16'h4472] = 8'hA9;
mem[16'h4473] = 8'h10;
mem[16'h4474] = 8'h20;
mem[16'h4475] = 8'h89;
mem[16'h4476] = 8'h66;
mem[16'h4477] = 8'hD8;
mem[16'h4478] = 8'h20;
mem[16'h4479] = 8'h0C;
mem[16'h447A] = 8'h4C;
mem[16'h447B] = 8'hF8;
mem[16'h447C] = 8'h4C;
mem[16'h447D] = 8'h66;
mem[16'h447E] = 8'h44;
mem[16'h447F] = 8'hD8;
mem[16'h4480] = 8'h20;
mem[16'h4481] = 8'h39;
mem[16'h4482] = 8'h49;
mem[16'h4483] = 8'h20;
mem[16'h4484] = 8'h97;
mem[16'h4485] = 8'h6E;
mem[16'h4486] = 8'hAD;
mem[16'h4487] = 8'h91;
mem[16'h4488] = 8'h6F;
mem[16'h4489] = 8'hF0;
mem[16'h448A] = 8'h0A;
mem[16'h448B] = 8'hA5;
mem[16'h448C] = 8'h60;
mem[16'h448D] = 8'hA4;
mem[16'h448E] = 8'h61;
mem[16'h448F] = 8'h20;
mem[16'h4490] = 8'h86;
mem[16'h4491] = 8'h68;
mem[16'h4492] = 8'h20;
mem[16'h4493] = 8'h37;
mem[16'h4494] = 8'h6F;
mem[16'h4495] = 8'hAD;
mem[16'h4496] = 8'hA8;
mem[16'h4497] = 8'h44;
mem[16'h4498] = 8'hC9;
mem[16'h4499] = 8'h05;
mem[16'h449A] = 8'hF0;
mem[16'h449B] = 8'h0E;
mem[16'h449C] = 8'h20;
mem[16'h449D] = 8'hFF;
mem[16'h449E] = 8'h44;
mem[16'h449F] = 8'h20;
mem[16'h44A0] = 8'hB4;
mem[16'h44A1] = 8'h4D;
mem[16'h44A2] = 8'h60;
mem[16'h44A3] = 8'h46;
mem[16'h44A4] = 8'hCB;
mem[16'h44A5] = 8'h15;
mem[16'h44A6] = 8'hA1;
mem[16'h44A7] = 8'h70;
mem[16'h44A8] = 8'h00;
mem[16'h44A9] = 8'h00;
mem[16'h44AA] = 8'h20;
mem[16'h44AB] = 8'hBE;
mem[16'h44AC] = 8'h41;
mem[16'h44AD] = 8'hA9;
mem[16'h44AE] = 8'h10;
mem[16'h44AF] = 8'h20;
mem[16'h44B0] = 8'hAD;
mem[16'h44B1] = 8'h66;
mem[16'h44B2] = 8'hEE;
mem[16'h44B3] = 8'hCE;
mem[16'h44B4] = 8'h44;
mem[16'h44B5] = 8'hAD;
mem[16'h44B6] = 8'hCE;
mem[16'h44B7] = 8'h44;
mem[16'h44B8] = 8'hA9;
mem[16'h44B9] = 8'hBA;
mem[16'h44BA] = 8'h85;
mem[16'h44BB] = 8'h79;
mem[16'h44BC] = 8'hA9;
mem[16'h44BD] = 8'h83;
mem[16'h44BE] = 8'h85;
mem[16'h44BF] = 8'h7A;
mem[16'h44C0] = 8'hA9;
mem[16'h44C1] = 8'hFB;
mem[16'h44C2] = 8'h85;
mem[16'h44C3] = 8'h7B;
mem[16'h44C4] = 8'hA9;
mem[16'h44C5] = 8'h83;
mem[16'h44C6] = 8'h85;
mem[16'h44C7] = 8'h7C;
mem[16'h44C8] = 8'h20;
mem[16'h44C9] = 8'hA2;
mem[16'h44CA] = 8'h82;
mem[16'h44CB] = 8'h4C;
mem[16'h44CC] = 8'h0F;
mem[16'h44CD] = 8'h40;
mem[16'h44CE] = 8'h01;
mem[16'h44CF] = 8'hA2;
mem[16'h44D0] = 8'h05;
mem[16'h44D1] = 8'hCA;
mem[16'h44D2] = 8'h30;
mem[16'h44D3] = 8'h2A;
mem[16'h44D4] = 8'hBD;
mem[16'h44D5] = 8'h5E;
mem[16'h44D6] = 8'h42;
mem[16'h44D7] = 8'hF0;
mem[16'h44D8] = 8'hF8;
mem[16'h44D9] = 8'hC9;
mem[16'h44DA] = 8'h01;
mem[16'h44DB] = 8'hF0;
mem[16'h44DC] = 8'h08;
mem[16'h44DD] = 8'hA9;
mem[16'h44DE] = 8'h00;
mem[16'h44DF] = 8'h9D;
mem[16'h44E0] = 8'h5E;
mem[16'h44E1] = 8'h42;
mem[16'h44E2] = 8'h4C;
mem[16'h44E3] = 8'hD1;
mem[16'h44E4] = 8'h44;
mem[16'h44E5] = 8'h86;
mem[16'h44E6] = 8'h70;
mem[16'h44E7] = 8'hA9;
mem[16'h44E8] = 8'h07;
mem[16'h44E9] = 8'h8D;
mem[16'h44EA] = 8'hD0;
mem[16'h44EB] = 8'h4D;
mem[16'h44EC] = 8'hBD;
mem[16'h44ED] = 8'hA3;
mem[16'h44EE] = 8'h44;
mem[16'h44EF] = 8'h8D;
mem[16'h44F0] = 8'hCF;
mem[16'h44F1] = 8'h4D;
mem[16'h44F2] = 8'hA9;
mem[16'h44F3] = 8'h00;
mem[16'h44F4] = 8'h85;
mem[16'h44F5] = 8'h77;
mem[16'h44F6] = 8'h20;
mem[16'h44F7] = 8'hD9;
mem[16'h44F8] = 8'h4C;
mem[16'h44F9] = 8'hA6;
mem[16'h44FA] = 8'h70;
mem[16'h44FB] = 8'h4C;
mem[16'h44FC] = 8'hD1;
mem[16'h44FD] = 8'h44;
mem[16'h44FE] = 8'h60;
mem[16'h44FF] = 8'hA9;
mem[16'h4500] = 8'h60;
mem[16'h4501] = 8'h85;
mem[16'h4502] = 8'h74;
mem[16'h4503] = 8'hA9;
mem[16'h4504] = 8'h05;
mem[16'h4505] = 8'h85;
mem[16'h4506] = 8'h73;
mem[16'h4507] = 8'hAD;
mem[16'h4508] = 8'hDF;
mem[16'h4509] = 8'h91;
mem[16'h450A] = 8'h8D;
mem[16'h450B] = 8'hDB;
mem[16'h450C] = 8'h91;
mem[16'h450D] = 8'hAD;
mem[16'h450E] = 8'hDD;
mem[16'h450F] = 8'h91;
mem[16'h4510] = 8'h8D;
mem[16'h4511] = 8'hDC;
mem[16'h4512] = 8'h91;
mem[16'h4513] = 8'hAD;
mem[16'h4514] = 8'hDE;
mem[16'h4515] = 8'h91;
mem[16'h4516] = 8'h8D;
mem[16'h4517] = 8'hDA;
mem[16'h4518] = 8'h91;
mem[16'h4519] = 8'hA0;
mem[16'h451A] = 8'h27;
mem[16'h451B] = 8'hA2;
mem[16'h451C] = 8'h46;
mem[16'h451D] = 8'h8E;
mem[16'h451E] = 8'h34;
mem[16'h451F] = 8'h45;
mem[16'h4520] = 8'hBD;
mem[16'h4521] = 8'hD5;
mem[16'h4522] = 8'h8E;
mem[16'h4523] = 8'h85;
mem[16'h4524] = 8'h59;
mem[16'h4525] = 8'hBD;
mem[16'h4526] = 8'h95;
mem[16'h4527] = 8'h8F;
mem[16'h4528] = 8'h85;
mem[16'h4529] = 8'h5A;
mem[16'h452A] = 8'hA9;
mem[16'h452B] = 8'h2A;
mem[16'h452C] = 8'h91;
mem[16'h452D] = 8'h59;
mem[16'h452E] = 8'hE8;
mem[16'h452F] = 8'hE0;
mem[16'h4530] = 8'hBE;
mem[16'h4531] = 8'hD0;
mem[16'h4532] = 8'hED;
mem[16'h4533] = 8'h60;
mem[16'h4534] = 8'h46;
mem[16'h4535] = 8'hAD;
mem[16'h4536] = 8'hD0;
mem[16'h4537] = 8'h4D;
mem[16'h4538] = 8'hC9;
mem[16'h4539] = 8'h4D;
mem[16'h453A] = 8'hD0;
mem[16'h453B] = 8'h44;
mem[16'h453C] = 8'hAE;
mem[16'h453D] = 8'hB0;
mem[16'h453E] = 8'h4A;
mem[16'h453F] = 8'hCA;
mem[16'h4540] = 8'hE0;
mem[16'h4541] = 8'h08;
mem[16'h4542] = 8'hB0;
mem[16'h4543] = 8'h03;
mem[16'h4544] = 8'h4C;
mem[16'h4545] = 8'h59;
mem[16'h4546] = 8'h48;
mem[16'h4547] = 8'hBD;
mem[16'h4548] = 8'h2C;
mem[16'h4549] = 8'h5F;
mem[16'h454A] = 8'h38;
mem[16'h454B] = 8'hE9;
mem[16'h454C] = 8'h0A;
mem[16'h454D] = 8'hB0;
mem[16'h454E] = 8'h02;
mem[16'h454F] = 8'hA9;
mem[16'h4550] = 8'h00;
mem[16'h4551] = 8'hCD;
mem[16'h4552] = 8'hCF;
mem[16'h4553] = 8'h4D;
mem[16'h4554] = 8'hB0;
mem[16'h4555] = 8'hE9;
mem[16'h4556] = 8'hBD;
mem[16'h4557] = 8'h2C;
mem[16'h4558] = 8'h5F;
mem[16'h4559] = 8'h18;
mem[16'h455A] = 8'h69;
mem[16'h455B] = 8'h10;
mem[16'h455C] = 8'h90;
mem[16'h455D] = 8'h02;
mem[16'h455E] = 8'hA9;
mem[16'h455F] = 8'hFF;
mem[16'h4560] = 8'hCD;
mem[16'h4561] = 8'hCF;
mem[16'h4562] = 8'h4D;
mem[16'h4563] = 8'h90;
mem[16'h4564] = 8'hDA;
mem[16'h4565] = 8'hBD;
mem[16'h4566] = 8'h75;
mem[16'h4567] = 8'h5B;
mem[16'h4568] = 8'hC9;
mem[16'h4569] = 8'h16;
mem[16'h456A] = 8'hB0;
mem[16'h456B] = 8'h07;
mem[16'h456C] = 8'hC9;
mem[16'h456D] = 8'h0F;
mem[16'h456E] = 8'h90;
mem[16'h456F] = 8'h03;
mem[16'h4570] = 8'h4C;
mem[16'h4571] = 8'h59;
mem[16'h4572] = 8'h48;
mem[16'h4573] = 8'hAD;
mem[16'h4574] = 8'hB6;
mem[16'h4575] = 8'h4A;
mem[16'h4576] = 8'hC9;
mem[16'h4577] = 8'h01;
mem[16'h4578] = 8'hD0;
mem[16'h4579] = 8'h03;
mem[16'h457A] = 8'h4C;
mem[16'h457B] = 8'hFE;
mem[16'h457C] = 8'h46;
mem[16'h457D] = 8'h4C;
mem[16'h457E] = 8'h14;
mem[16'h457F] = 8'h47;
mem[16'h4580] = 8'hC9;
mem[16'h4581] = 8'h23;
mem[16'h4582] = 8'hD0;
mem[16'h4583] = 8'h49;
mem[16'h4584] = 8'hAE;
mem[16'h4585] = 8'hAF;
mem[16'h4586] = 8'h4A;
mem[16'h4587] = 8'hCA;
mem[16'h4588] = 8'h30;
mem[16'h4589] = 8'h40;
mem[16'h458A] = 8'hBD;
mem[16'h458B] = 8'h2C;
mem[16'h458C] = 8'h5F;
mem[16'h458D] = 8'h38;
mem[16'h458E] = 8'hE9;
mem[16'h458F] = 8'h0A;
mem[16'h4590] = 8'hB0;
mem[16'h4591] = 8'h02;
mem[16'h4592] = 8'hA9;
mem[16'h4593] = 8'h00;
mem[16'h4594] = 8'hCD;
mem[16'h4595] = 8'hCF;
mem[16'h4596] = 8'h4D;
mem[16'h4597] = 8'hB0;
mem[16'h4598] = 8'hEE;
mem[16'h4599] = 8'hBD;
mem[16'h459A] = 8'h2C;
mem[16'h459B] = 8'h5F;
mem[16'h459C] = 8'h18;
mem[16'h459D] = 8'h69;
mem[16'h459E] = 8'h10;
mem[16'h459F] = 8'h90;
mem[16'h45A0] = 8'h02;
mem[16'h45A1] = 8'hA9;
mem[16'h45A2] = 8'hFF;
mem[16'h45A3] = 8'hCD;
mem[16'h45A4] = 8'hCF;
mem[16'h45A5] = 8'h4D;
mem[16'h45A6] = 8'h90;
mem[16'h45A7] = 8'hDF;
mem[16'h45A8] = 8'hBD;
mem[16'h45A9] = 8'h75;
mem[16'h45AA] = 8'h5B;
mem[16'h45AB] = 8'hC9;
mem[16'h45AC] = 8'h16;
mem[16'h45AD] = 8'hB0;
mem[16'h45AE] = 8'h07;
mem[16'h45AF] = 8'hC9;
mem[16'h45B0] = 8'h0F;
mem[16'h45B1] = 8'h90;
mem[16'h45B2] = 8'h03;
mem[16'h45B3] = 8'h4C;
mem[16'h45B4] = 8'h59;
mem[16'h45B5] = 8'h48;
mem[16'h45B6] = 8'hAD;
mem[16'h45B7] = 8'hB7;
mem[16'h45B8] = 8'h4A;
mem[16'h45B9] = 8'hC9;
mem[16'h45BA] = 8'h01;
mem[16'h45BB] = 8'hD0;
mem[16'h45BC] = 8'h09;
mem[16'h45BD] = 8'hA5;
mem[16'h45BE] = 8'h73;
mem[16'h45BF] = 8'h29;
mem[16'h45C0] = 8'h01;
mem[16'h45C1] = 8'hF0;
mem[16'h45C2] = 8'h03;
mem[16'h45C3] = 8'h4C;
mem[16'h45C4] = 8'hFE;
mem[16'h45C5] = 8'h46;
mem[16'h45C6] = 8'h4C;
mem[16'h45C7] = 8'h14;
mem[16'h45C8] = 8'h47;
mem[16'h45C9] = 8'h60;
mem[16'h45CA] = 8'h4C;
mem[16'h45CB] = 8'h59;
mem[16'h45CC] = 8'h48;
mem[16'h45CD] = 8'hC9;
mem[16'h45CE] = 8'h3F;
mem[16'h45CF] = 8'hD0;
mem[16'h45D0] = 8'h2B;
mem[16'h45D1] = 8'hAE;
mem[16'h45D2] = 8'hB3;
mem[16'h45D3] = 8'h4A;
mem[16'h45D4] = 8'hCA;
mem[16'h45D5] = 8'h30;
mem[16'h45D6] = 8'hF3;
mem[16'h45D7] = 8'hBD;
mem[16'h45D8] = 8'h1F;
mem[16'h45D9] = 8'h53;
mem[16'h45DA] = 8'h38;
mem[16'h45DB] = 8'hE9;
mem[16'h45DC] = 8'h02;
mem[16'h45DD] = 8'hCD;
mem[16'h45DE] = 8'hCF;
mem[16'h45DF] = 8'h4D;
mem[16'h45E0] = 8'h90;
mem[16'h45E1] = 8'hF2;
mem[16'h45E2] = 8'hBD;
mem[16'h45E3] = 8'h1F;
mem[16'h45E4] = 8'h53;
mem[16'h45E5] = 8'h38;
mem[16'h45E6] = 8'hFD;
mem[16'h45E7] = 8'h28;
mem[16'h45E8] = 8'h53;
mem[16'h45E9] = 8'h90;
mem[16'h45EA] = 8'h07;
mem[16'h45EB] = 8'hE9;
mem[16'h45EC] = 8'h0B;
mem[16'h45ED] = 8'h90;
mem[16'h45EE] = 8'h03;
mem[16'h45EF] = 8'h4C;
mem[16'h45F0] = 8'hF4;
mem[16'h45F1] = 8'h45;
mem[16'h45F2] = 8'hA9;
mem[16'h45F3] = 8'h00;
mem[16'h45F4] = 8'hCD;
mem[16'h45F5] = 8'hCF;
mem[16'h45F6] = 8'h4D;
mem[16'h45F7] = 8'hB0;
mem[16'h45F8] = 8'hDB;
mem[16'h45F9] = 8'h4C;
mem[16'h45FA] = 8'hC8;
mem[16'h45FB] = 8'h46;
mem[16'h45FC] = 8'hC9;
mem[16'h45FD] = 8'h31;
mem[16'h45FE] = 8'hD0;
mem[16'h45FF] = 8'h4B;
mem[16'h4600] = 8'hAE;
mem[16'h4601] = 8'hB2;
mem[16'h4602] = 8'h4A;
mem[16'h4603] = 8'hCA;
mem[16'h4604] = 8'h30;
mem[16'h4605] = 8'hC4;
mem[16'h4606] = 8'hBD;
mem[16'h4607] = 8'h10;
mem[16'h4608] = 8'h51;
mem[16'h4609] = 8'h38;
mem[16'h460A] = 8'hE9;
mem[16'h460B] = 8'h02;
mem[16'h460C] = 8'hCD;
mem[16'h460D] = 8'hCF;
mem[16'h460E] = 8'h4D;
mem[16'h460F] = 8'h90;
mem[16'h4610] = 8'h24;
mem[16'h4611] = 8'hBD;
mem[16'h4612] = 8'h10;
mem[16'h4613] = 8'h51;
mem[16'h4614] = 8'h38;
mem[16'h4615] = 8'hFD;
mem[16'h4616] = 8'h16;
mem[16'h4617] = 8'h51;
mem[16'h4618] = 8'h90;
mem[16'h4619] = 8'h07;
mem[16'h461A] = 8'hE9;
mem[16'h461B] = 8'h0B;
mem[16'h461C] = 8'h90;
mem[16'h461D] = 8'h03;
mem[16'h461E] = 8'h4C;
mem[16'h461F] = 8'h23;
mem[16'h4620] = 8'h46;
mem[16'h4621] = 8'hA9;
mem[16'h4622] = 8'h00;
mem[16'h4623] = 8'hCD;
mem[16'h4624] = 8'hCF;
mem[16'h4625] = 8'h4D;
mem[16'h4626] = 8'hB0;
mem[16'h4627] = 8'hDB;
mem[16'h4628] = 8'hAD;
mem[16'h4629] = 8'hB5;
mem[16'h462A] = 8'h4A;
mem[16'h462B] = 8'hC9;
mem[16'h462C] = 8'h01;
mem[16'h462D] = 8'hD0;
mem[16'h462E] = 8'h03;
mem[16'h462F] = 8'h4C;
mem[16'h4630] = 8'hE3;
mem[16'h4631] = 8'h46;
mem[16'h4632] = 8'h4C;
mem[16'h4633] = 8'h2A;
mem[16'h4634] = 8'h47;
mem[16'h4635] = 8'hAC;
mem[16'h4636] = 8'hB2;
mem[16'h4637] = 8'h4A;
mem[16'h4638] = 8'hC0;
mem[16'h4639] = 8'h01;
mem[16'h463A] = 8'hD0;
mem[16'h463B] = 8'hC7;
mem[16'h463C] = 8'hBD;
mem[16'h463D] = 8'h10;
mem[16'h463E] = 8'h51;
mem[16'h463F] = 8'h38;
mem[16'h4640] = 8'hFD;
mem[16'h4641] = 8'h16;
mem[16'h4642] = 8'h51;
mem[16'h4643] = 8'hB0;
mem[16'h4644] = 8'hBE;
mem[16'h4645] = 8'h38;
mem[16'h4646] = 8'hE9;
mem[16'h4647] = 8'h0B;
mem[16'h4648] = 8'h4C;
mem[16'h4649] = 8'h23;
mem[16'h464A] = 8'h46;
mem[16'h464B] = 8'hC9;
mem[16'h464C] = 8'h15;
mem[16'h464D] = 8'hD0;
mem[16'h464E] = 8'h65;
mem[16'h464F] = 8'hAE;
mem[16'h4650] = 8'hB1;
mem[16'h4651] = 8'h4A;
mem[16'h4652] = 8'hCA;
mem[16'h4653] = 8'h30;
mem[16'h4654] = 8'h35;
mem[16'h4655] = 8'hBD;
mem[16'h4656] = 8'h00;
mem[16'h4657] = 8'h54;
mem[16'h4658] = 8'h38;
mem[16'h4659] = 8'hE9;
mem[16'h465A] = 8'h02;
mem[16'h465B] = 8'hCD;
mem[16'h465C] = 8'hCF;
mem[16'h465D] = 8'h4D;
mem[16'h465E] = 8'h90;
mem[16'h465F] = 8'hF2;
mem[16'h4660] = 8'hBD;
mem[16'h4661] = 8'h00;
mem[16'h4662] = 8'h54;
mem[16'h4663] = 8'h38;
mem[16'h4664] = 8'hFD;
mem[16'h4665] = 8'h0D;
mem[16'h4666] = 8'h54;
mem[16'h4667] = 8'h90;
mem[16'h4668] = 8'h07;
mem[16'h4669] = 8'hE9;
mem[16'h466A] = 8'h0B;
mem[16'h466B] = 8'h90;
mem[16'h466C] = 8'h03;
mem[16'h466D] = 8'h4C;
mem[16'h466E] = 8'h72;
mem[16'h466F] = 8'h46;
mem[16'h4670] = 8'hA9;
mem[16'h4671] = 8'h00;
mem[16'h4672] = 8'hCD;
mem[16'h4673] = 8'hCF;
mem[16'h4674] = 8'h4D;
mem[16'h4675] = 8'hB0;
mem[16'h4676] = 8'hDB;
mem[16'h4677] = 8'hAD;
mem[16'h4678] = 8'hB4;
mem[16'h4679] = 8'h4A;
mem[16'h467A] = 8'hC9;
mem[16'h467B] = 8'h01;
mem[16'h467C] = 8'hF0;
mem[16'h467D] = 8'h09;
mem[16'h467E] = 8'hA5;
mem[16'h467F] = 8'h73;
mem[16'h4680] = 8'h29;
mem[16'h4681] = 8'h01;
mem[16'h4682] = 8'hD0;
mem[16'h4683] = 8'h03;
mem[16'h4684] = 8'h4C;
mem[16'h4685] = 8'hE3;
mem[16'h4686] = 8'h46;
mem[16'h4687] = 8'h4C;
mem[16'h4688] = 8'hC8;
mem[16'h4689] = 8'h46;
mem[16'h468A] = 8'hAE;
mem[16'h468B] = 8'h5A;
mem[16'h468C] = 8'h74;
mem[16'h468D] = 8'hCA;
mem[16'h468E] = 8'h30;
mem[16'h468F] = 8'h25;
mem[16'h4690] = 8'hBD;
mem[16'h4691] = 8'h84;
mem[16'h4692] = 8'h7B;
mem[16'h4693] = 8'h38;
mem[16'h4694] = 8'hE9;
mem[16'h4695] = 8'h0A;
mem[16'h4696] = 8'hCD;
mem[16'h4697] = 8'hCF;
mem[16'h4698] = 8'h4D;
mem[16'h4699] = 8'hB0;
mem[16'h469A] = 8'hF2;
mem[16'h469B] = 8'hBD;
mem[16'h469C] = 8'h84;
mem[16'h469D] = 8'h7B;
mem[16'h469E] = 8'h18;
mem[16'h469F] = 8'h69;
mem[16'h46A0] = 8'h18;
mem[16'h46A1] = 8'hCD;
mem[16'h46A2] = 8'hCF;
mem[16'h46A3] = 8'h4D;
mem[16'h46A4] = 8'hB0;
mem[16'h46A5] = 8'h12;
mem[16'h46A6] = 8'hBD;
mem[16'h46A7] = 8'h84;
mem[16'h46A8] = 8'h7B;
mem[16'h46A9] = 8'h18;
mem[16'h46AA] = 8'h69;
mem[16'h46AB] = 8'h31;
mem[16'h46AC] = 8'hCD;
mem[16'h46AD] = 8'hCF;
mem[16'h46AE] = 8'h4D;
mem[16'h46AF] = 8'h90;
mem[16'h46B0] = 8'hDC;
mem[16'h46B1] = 8'h4C;
mem[16'h46B2] = 8'h8E;
mem[16'h46B3] = 8'h48;
mem[16'h46B4] = 8'h60;
mem[16'h46B5] = 8'h4C;
mem[16'h46B6] = 8'h59;
mem[16'h46B7] = 8'h48;
mem[16'h46B8] = 8'hAD;
mem[16'h46B9] = 8'hB4;
mem[16'h46BA] = 8'h4A;
mem[16'h46BB] = 8'hC9;
mem[16'h46BC] = 8'h01;
mem[16'h46BD] = 8'hF0;
mem[16'h46BE] = 8'h09;
mem[16'h46BF] = 8'hA5;
mem[16'h46C0] = 8'h73;
mem[16'h46C1] = 8'h29;
mem[16'h46C2] = 8'h01;
mem[16'h46C3] = 8'hD0;
mem[16'h46C4] = 8'h03;
mem[16'h46C5] = 8'h4C;
mem[16'h46C6] = 8'hE3;
mem[16'h46C7] = 8'h46;
mem[16'h46C8] = 8'hAD;
mem[16'h46C9] = 8'hCF;
mem[16'h46CA] = 8'h4D;
mem[16'h46CB] = 8'hC9;
mem[16'h46CC] = 8'hFF;
mem[16'h46CD] = 8'hF0;
mem[16'h46CE] = 8'hE6;
mem[16'h46CF] = 8'h20;
mem[16'h46D0] = 8'hAE;
mem[16'h46D1] = 8'h4C;
mem[16'h46D2] = 8'hAD;
mem[16'h46D3] = 8'hCF;
mem[16'h46D4] = 8'h4D;
mem[16'h46D5] = 8'h18;
mem[16'h46D6] = 8'h69;
mem[16'h46D7] = 8'h02;
mem[16'h46D8] = 8'h90;
mem[16'h46D9] = 8'h02;
mem[16'h46DA] = 8'hA9;
mem[16'h46DB] = 8'hFF;
mem[16'h46DC] = 8'h8D;
mem[16'h46DD] = 8'hCF;
mem[16'h46DE] = 8'h4D;
mem[16'h46DF] = 8'h20;
mem[16'h46E0] = 8'hAE;
mem[16'h46E1] = 8'h4C;
mem[16'h46E2] = 8'h60;
mem[16'h46E3] = 8'hAD;
mem[16'h46E4] = 8'hCF;
mem[16'h46E5] = 8'h4D;
mem[16'h46E6] = 8'hC9;
mem[16'h46E7] = 8'hFF;
mem[16'h46E8] = 8'hF0;
mem[16'h46E9] = 8'hCB;
mem[16'h46EA] = 8'h20;
mem[16'h46EB] = 8'hAE;
mem[16'h46EC] = 8'h4C;
mem[16'h46ED] = 8'hAD;
mem[16'h46EE] = 8'hCF;
mem[16'h46EF] = 8'h4D;
mem[16'h46F0] = 8'h18;
mem[16'h46F1] = 8'h69;
mem[16'h46F2] = 8'h04;
mem[16'h46F3] = 8'h90;
mem[16'h46F4] = 8'h02;
mem[16'h46F5] = 8'hA9;
mem[16'h46F6] = 8'hFF;
mem[16'h46F7] = 8'h8D;
mem[16'h46F8] = 8'hCF;
mem[16'h46F9] = 8'h4D;
mem[16'h46FA] = 8'h20;
mem[16'h46FB] = 8'hAE;
mem[16'h46FC] = 8'h4C;
mem[16'h46FD] = 8'h60;
mem[16'h46FE] = 8'h20;
mem[16'h46FF] = 8'hAE;
mem[16'h4700] = 8'h4C;
mem[16'h4701] = 8'hAD;
mem[16'h4702] = 8'hCF;
mem[16'h4703] = 8'h4D;
mem[16'h4704] = 8'hF0;
mem[16'h4705] = 8'h07;
mem[16'h4706] = 8'h38;
mem[16'h4707] = 8'hE9;
mem[16'h4708] = 8'h02;
mem[16'h4709] = 8'hB0;
mem[16'h470A] = 8'h02;
mem[16'h470B] = 8'hA9;
mem[16'h470C] = 8'h00;
mem[16'h470D] = 8'h8D;
mem[16'h470E] = 8'hCF;
mem[16'h470F] = 8'h4D;
mem[16'h4710] = 8'h20;
mem[16'h4711] = 8'hAE;
mem[16'h4712] = 8'h4C;
mem[16'h4713] = 8'h60;
mem[16'h4714] = 8'h20;
mem[16'h4715] = 8'hAE;
mem[16'h4716] = 8'h4C;
mem[16'h4717] = 8'hAD;
mem[16'h4718] = 8'hCF;
mem[16'h4719] = 8'h4D;
mem[16'h471A] = 8'hF0;
mem[16'h471B] = 8'h07;
mem[16'h471C] = 8'h38;
mem[16'h471D] = 8'hE9;
mem[16'h471E] = 8'h04;
mem[16'h471F] = 8'hB0;
mem[16'h4720] = 8'h02;
mem[16'h4721] = 8'hA9;
mem[16'h4722] = 8'h00;
mem[16'h4723] = 8'h8D;
mem[16'h4724] = 8'hCF;
mem[16'h4725] = 8'h4D;
mem[16'h4726] = 8'h20;
mem[16'h4727] = 8'hAE;
mem[16'h4728] = 8'h4C;
mem[16'h4729] = 8'h60;
mem[16'h472A] = 8'hAD;
mem[16'h472B] = 8'hCF;
mem[16'h472C] = 8'h4D;
mem[16'h472D] = 8'hC9;
mem[16'h472E] = 8'hFF;
mem[16'h472F] = 8'hD0;
mem[16'h4730] = 8'h03;
mem[16'h4731] = 8'h4C;
mem[16'h4732] = 8'h59;
mem[16'h4733] = 8'h48;
mem[16'h4734] = 8'h20;
mem[16'h4735] = 8'hAE;
mem[16'h4736] = 8'h4C;
mem[16'h4737] = 8'hAD;
mem[16'h4738] = 8'hCF;
mem[16'h4739] = 8'h4D;
mem[16'h473A] = 8'h18;
mem[16'h473B] = 8'h69;
mem[16'h473C] = 8'h08;
mem[16'h473D] = 8'h90;
mem[16'h473E] = 8'h02;
mem[16'h473F] = 8'hA9;
mem[16'h4740] = 8'hFF;
mem[16'h4741] = 8'h8D;
mem[16'h4742] = 8'hCF;
mem[16'h4743] = 8'h4D;
mem[16'h4744] = 8'h20;
mem[16'h4745] = 8'hAE;
mem[16'h4746] = 8'h4C;
mem[16'h4747] = 8'h60;
mem[16'h4748] = 8'hAE;
mem[16'h4749] = 8'hAC;
mem[16'h474A] = 8'h4A;
mem[16'h474B] = 8'hCA;
mem[16'h474C] = 8'h30;
mem[16'h474D] = 8'h1F;
mem[16'h474E] = 8'hBD;
mem[16'h474F] = 8'h2E;
mem[16'h4750] = 8'h61;
mem[16'h4751] = 8'h38;
mem[16'h4752] = 8'hED;
mem[16'h4753] = 8'hD0;
mem[16'h4754] = 8'h4D;
mem[16'h4755] = 8'h20;
mem[16'h4756] = 8'h62;
mem[16'h4757] = 8'h65;
mem[16'h4758] = 8'hC9;
mem[16'h4759] = 8'h09;
mem[16'h475A] = 8'hB0;
mem[16'h475B] = 8'hEF;
mem[16'h475C] = 8'hBD;
mem[16'h475D] = 8'h2A;
mem[16'h475E] = 8'h61;
mem[16'h475F] = 8'h38;
mem[16'h4760] = 8'hED;
mem[16'h4761] = 8'hCF;
mem[16'h4762] = 8'h4D;
mem[16'h4763] = 8'h20;
mem[16'h4764] = 8'h62;
mem[16'h4765] = 8'h65;
mem[16'h4766] = 8'hC9;
mem[16'h4767] = 8'h0F;
mem[16'h4768] = 8'hB0;
mem[16'h4769] = 8'hE1;
mem[16'h476A] = 8'h4C;
mem[16'h476B] = 8'h79;
mem[16'h476C] = 8'h48;
mem[16'h476D] = 8'hAE;
mem[16'h476E] = 8'hAB;
mem[16'h476F] = 8'h4A;
mem[16'h4770] = 8'hCA;
mem[16'h4771] = 8'h30;
mem[16'h4772] = 8'h1F;
mem[16'h4773] = 8'hBD;
mem[16'h4774] = 8'hEF;
mem[16'h4775] = 8'h60;
mem[16'h4776] = 8'h38;
mem[16'h4777] = 8'hED;
mem[16'h4778] = 8'hD0;
mem[16'h4779] = 8'h4D;
mem[16'h477A] = 8'h20;
mem[16'h477B] = 8'h62;
mem[16'h477C] = 8'h65;
mem[16'h477D] = 8'hC9;
mem[16'h477E] = 8'h0A;
mem[16'h477F] = 8'hB0;
mem[16'h4780] = 8'hEF;
mem[16'h4781] = 8'hBD;
mem[16'h4782] = 8'hEB;
mem[16'h4783] = 8'h60;
mem[16'h4784] = 8'h38;
mem[16'h4785] = 8'hED;
mem[16'h4786] = 8'hCF;
mem[16'h4787] = 8'h4D;
mem[16'h4788] = 8'h20;
mem[16'h4789] = 8'h62;
mem[16'h478A] = 8'h65;
mem[16'h478B] = 8'hC9;
mem[16'h478C] = 8'h0F;
mem[16'h478D] = 8'hB0;
mem[16'h478E] = 8'hE1;
mem[16'h478F] = 8'h4C;
mem[16'h4790] = 8'h79;
mem[16'h4791] = 8'h48;
mem[16'h4792] = 8'hAE;
mem[16'h4793] = 8'hAA;
mem[16'h4794] = 8'h4A;
mem[16'h4795] = 8'hCA;
mem[16'h4796] = 8'h30;
mem[16'h4797] = 8'h1F;
mem[16'h4798] = 8'hBD;
mem[16'h4799] = 8'hAB;
mem[16'h479A] = 8'h60;
mem[16'h479B] = 8'h38;
mem[16'h479C] = 8'hED;
mem[16'h479D] = 8'hD0;
mem[16'h479E] = 8'h4D;
mem[16'h479F] = 8'h20;
mem[16'h47A0] = 8'h62;
mem[16'h47A1] = 8'h65;
mem[16'h47A2] = 8'hC9;
mem[16'h47A3] = 8'h0A;
mem[16'h47A4] = 8'hB0;
mem[16'h47A5] = 8'hEF;
mem[16'h47A6] = 8'hBD;
mem[16'h47A7] = 8'hA7;
mem[16'h47A8] = 8'h60;
mem[16'h47A9] = 8'h38;
mem[16'h47AA] = 8'hED;
mem[16'h47AB] = 8'hCF;
mem[16'h47AC] = 8'h4D;
mem[16'h47AD] = 8'h20;
mem[16'h47AE] = 8'h62;
mem[16'h47AF] = 8'h65;
mem[16'h47B0] = 8'hC9;
mem[16'h47B1] = 8'h0C;
mem[16'h47B2] = 8'hB0;
mem[16'h47B3] = 8'hE1;
mem[16'h47B4] = 8'h4C;
mem[16'h47B5] = 8'h79;
mem[16'h47B6] = 8'h48;
mem[16'h47B7] = 8'hAE;
mem[16'h47B8] = 8'hAD;
mem[16'h47B9] = 8'h4A;
mem[16'h47BA] = 8'hCA;
mem[16'h47BB] = 8'h30;
mem[16'h47BC] = 8'h1F;
mem[16'h47BD] = 8'hBD;
mem[16'h47BE] = 8'hB3;
mem[16'h47BF] = 8'h60;
mem[16'h47C0] = 8'h38;
mem[16'h47C1] = 8'hED;
mem[16'h47C2] = 8'hD0;
mem[16'h47C3] = 8'h4D;
mem[16'h47C4] = 8'h20;
mem[16'h47C5] = 8'h62;
mem[16'h47C6] = 8'h65;
mem[16'h47C7] = 8'hC9;
mem[16'h47C8] = 8'h0A;
mem[16'h47C9] = 8'hB0;
mem[16'h47CA] = 8'hEF;
mem[16'h47CB] = 8'hBD;
mem[16'h47CC] = 8'hAF;
mem[16'h47CD] = 8'h60;
mem[16'h47CE] = 8'h38;
mem[16'h47CF] = 8'hED;
mem[16'h47D0] = 8'hCF;
mem[16'h47D1] = 8'h4D;
mem[16'h47D2] = 8'h20;
mem[16'h47D3] = 8'h62;
mem[16'h47D4] = 8'h65;
mem[16'h47D5] = 8'hC9;
mem[16'h47D6] = 8'h0F;
mem[16'h47D7] = 8'hB0;
mem[16'h47D8] = 8'hE1;
mem[16'h47D9] = 8'h4C;
mem[16'h47DA] = 8'h79;
mem[16'h47DB] = 8'h48;
mem[16'h47DC] = 8'hAE;
mem[16'h47DD] = 8'hAE;
mem[16'h47DE] = 8'h4A;
mem[16'h47DF] = 8'hCA;
mem[16'h47E0] = 8'h30;
mem[16'h47E1] = 8'h1F;
mem[16'h47E2] = 8'hBD;
mem[16'h47E3] = 8'h4A;
mem[16'h47E4] = 8'h60;
mem[16'h47E5] = 8'h38;
mem[16'h47E6] = 8'hED;
mem[16'h47E7] = 8'hD0;
mem[16'h47E8] = 8'h4D;
mem[16'h47E9] = 8'h20;
mem[16'h47EA] = 8'h62;
mem[16'h47EB] = 8'h65;
mem[16'h47EC] = 8'hC9;
mem[16'h47ED] = 8'h0A;
mem[16'h47EE] = 8'hB0;
mem[16'h47EF] = 8'hEF;
mem[16'h47F0] = 8'hBD;
mem[16'h47F1] = 8'h47;
mem[16'h47F2] = 8'h60;
mem[16'h47F3] = 8'h38;
mem[16'h47F4] = 8'hED;
mem[16'h47F5] = 8'hCF;
mem[16'h47F6] = 8'h4D;
mem[16'h47F7] = 8'h20;
mem[16'h47F8] = 8'h62;
mem[16'h47F9] = 8'h65;
mem[16'h47FA] = 8'hC9;
mem[16'h47FB] = 8'h0F;
mem[16'h47FC] = 8'hB0;
mem[16'h47FD] = 8'hE1;
mem[16'h47FE] = 8'h4C;
mem[16'h47FF] = 8'h79;
mem[16'h4800] = 8'h48;
mem[16'h4801] = 8'hAD;
mem[16'h4802] = 8'hC0;
mem[16'h4803] = 8'h62;
mem[16'h4804] = 8'hF0;
mem[16'h4805] = 8'h24;
mem[16'h4806] = 8'hAD;
mem[16'h4807] = 8'hBA;
mem[16'h4808] = 8'h62;
mem[16'h4809] = 8'h38;
mem[16'h480A] = 8'hED;
mem[16'h480B] = 8'hD0;
mem[16'h480C] = 8'h4D;
mem[16'h480D] = 8'h20;
mem[16'h480E] = 8'h62;
mem[16'h480F] = 8'h65;
mem[16'h4810] = 8'hC9;
mem[16'h4811] = 8'h05;
mem[16'h4812] = 8'hB0;
mem[16'h4813] = 8'h16;
mem[16'h4814] = 8'hAD;
mem[16'h4815] = 8'hB8;
mem[16'h4816] = 8'h62;
mem[16'h4817] = 8'h18;
mem[16'h4818] = 8'h69;
mem[16'h4819] = 8'h01;
mem[16'h481A] = 8'hCD;
mem[16'h481B] = 8'hCF;
mem[16'h481C] = 8'h4D;
mem[16'h481D] = 8'hB0;
mem[16'h481E] = 8'h0B;
mem[16'h481F] = 8'h18;
mem[16'h4820] = 8'h69;
mem[16'h4821] = 8'h15;
mem[16'h4822] = 8'hCD;
mem[16'h4823] = 8'hCF;
mem[16'h4824] = 8'h4D;
mem[16'h4825] = 8'h90;
mem[16'h4826] = 8'h03;
mem[16'h4827] = 8'h4C;
mem[16'h4828] = 8'h8E;
mem[16'h4829] = 8'h48;
mem[16'h482A] = 8'hA2;
mem[16'h482B] = 8'h02;
mem[16'h482C] = 8'hCA;
mem[16'h482D] = 8'h30;
mem[16'h482E] = 8'h29;
mem[16'h482F] = 8'hBD;
mem[16'h4830] = 8'hC2;
mem[16'h4831] = 8'h62;
mem[16'h4832] = 8'hF0;
mem[16'h4833] = 8'hF8;
mem[16'h4834] = 8'hBD;
mem[16'h4835] = 8'hBE;
mem[16'h4836] = 8'h62;
mem[16'h4837] = 8'h38;
mem[16'h4838] = 8'hED;
mem[16'h4839] = 8'hD0;
mem[16'h483A] = 8'h4D;
mem[16'h483B] = 8'h20;
mem[16'h483C] = 8'h62;
mem[16'h483D] = 8'h65;
mem[16'h483E] = 8'hC9;
mem[16'h483F] = 8'h05;
mem[16'h4840] = 8'hB0;
mem[16'h4841] = 8'hEA;
mem[16'h4842] = 8'hBD;
mem[16'h4843] = 8'hBC;
mem[16'h4844] = 8'h62;
mem[16'h4845] = 8'h18;
mem[16'h4846] = 8'h69;
mem[16'h4847] = 8'h07;
mem[16'h4848] = 8'hCD;
mem[16'h4849] = 8'hCF;
mem[16'h484A] = 8'h4D;
mem[16'h484B] = 8'h90;
mem[16'h484C] = 8'hDF;
mem[16'h484D] = 8'h38;
mem[16'h484E] = 8'hE9;
mem[16'h484F] = 8'h13;
mem[16'h4850] = 8'hCD;
mem[16'h4851] = 8'hCF;
mem[16'h4852] = 8'h4D;
mem[16'h4853] = 8'hB0;
mem[16'h4854] = 8'hD7;
mem[16'h4855] = 8'h4C;
mem[16'h4856] = 8'h8E;
mem[16'h4857] = 8'h48;
mem[16'h4858] = 8'h60;
mem[16'h4859] = 8'hA9;
mem[16'h485A] = 8'h00;
mem[16'h485B] = 8'h8D;
mem[16'h485C] = 8'h2E;
mem[16'h485D] = 8'h49;
mem[16'h485E] = 8'h20;
mem[16'h485F] = 8'hAE;
mem[16'h4860] = 8'h4C;
mem[16'h4861] = 8'h20;
mem[16'h4862] = 8'hEF;
mem[16'h4863] = 8'h4B;
mem[16'h4864] = 8'h20;
mem[16'h4865] = 8'h01;
mem[16'h4866] = 8'h49;
mem[16'h4867] = 8'h20;
mem[16'h4868] = 8'h01;
mem[16'h4869] = 8'h49;
mem[16'h486A] = 8'h20;
mem[16'h486B] = 8'h01;
mem[16'h486C] = 8'h49;
mem[16'h486D] = 8'h20;
mem[16'h486E] = 8'h01;
mem[16'h486F] = 8'h49;
mem[16'h4870] = 8'h20;
mem[16'h4871] = 8'h01;
mem[16'h4872] = 8'h49;
mem[16'h4873] = 8'h20;
mem[16'h4874] = 8'hBE;
mem[16'h4875] = 8'h7E;
mem[16'h4876] = 8'h4C;
mem[16'h4877] = 8'h97;
mem[16'h4878] = 8'h48;
mem[16'h4879] = 8'h20;
mem[16'h487A] = 8'hAE;
mem[16'h487B] = 8'h4C;
mem[16'h487C] = 8'h20;
mem[16'h487D] = 8'hE7;
mem[16'h487E] = 8'h48;
mem[16'h487F] = 8'h20;
mem[16'h4880] = 8'h4A;
mem[16'h4881] = 8'h4C;
mem[16'h4882] = 8'h20;
mem[16'h4883] = 8'h47;
mem[16'h4884] = 8'h49;
mem[16'h4885] = 8'h20;
mem[16'h4886] = 8'hE7;
mem[16'h4887] = 8'h48;
mem[16'h4888] = 8'h20;
mem[16'h4889] = 8'hBE;
mem[16'h488A] = 8'h7E;
mem[16'h488B] = 8'h4C;
mem[16'h488C] = 8'h97;
mem[16'h488D] = 8'h48;
mem[16'h488E] = 8'h20;
mem[16'h488F] = 8'hAE;
mem[16'h4890] = 8'h4C;
mem[16'h4891] = 8'h20;
mem[16'h4892] = 8'hBE;
mem[16'h4893] = 8'h7E;
mem[16'h4894] = 8'h20;
mem[16'h4895] = 8'h6D;
mem[16'h4896] = 8'h4C;
mem[16'h4897] = 8'h20;
mem[16'h4898] = 8'h39;
mem[16'h4899] = 8'h49;
mem[16'h489A] = 8'hAD;
mem[16'h489B] = 8'hB3;
mem[16'h489C] = 8'h85;
mem[16'h489D] = 8'hF0;
mem[16'h489E] = 8'h08;
mem[16'h489F] = 8'h20;
mem[16'h48A0] = 8'h0E;
mem[16'h48A1] = 8'h73;
mem[16'h48A2] = 8'hA9;
mem[16'h48A3] = 8'h00;
mem[16'h48A4] = 8'h8D;
mem[16'h48A5] = 8'hB3;
mem[16'h48A6] = 8'h85;
mem[16'h48A7] = 8'hCE;
mem[16'h48A8] = 8'hE6;
mem[16'h48A9] = 8'h48;
mem[16'h48AA] = 8'hF0;
mem[16'h48AB] = 8'h2D;
mem[16'h48AC] = 8'hA5;
mem[16'h48AD] = 8'h74;
mem[16'h48AE] = 8'hD0;
mem[16'h48AF] = 8'h06;
mem[16'h48B0] = 8'h20;
mem[16'h48B1] = 8'hED;
mem[16'h48B2] = 8'h6D;
mem[16'h48B3] = 8'h4C;
mem[16'h48B4] = 8'hB9;
mem[16'h48B5] = 8'h48;
mem[16'h48B6] = 8'h20;
mem[16'h48B7] = 8'hBE;
mem[16'h48B8] = 8'h7E;
mem[16'h48B9] = 8'h20;
mem[16'h48BA] = 8'hFF;
mem[16'h48BB] = 8'h44;
mem[16'h48BC] = 8'hAD;
mem[16'h48BD] = 8'hD3;
mem[16'h48BE] = 8'h90;
mem[16'h48BF] = 8'h85;
mem[16'h48C0] = 8'h56;
mem[16'h48C1] = 8'h38;
mem[16'h48C2] = 8'hE9;
mem[16'h48C3] = 8'h0E;
mem[16'h48C4] = 8'h8D;
mem[16'h48C5] = 8'hD3;
mem[16'h48C6] = 8'h90;
mem[16'h48C7] = 8'h20;
mem[16'h48C8] = 8'h54;
mem[16'h48C9] = 8'h8B;
mem[16'h48CA] = 8'h20;
mem[16'h48CB] = 8'hB4;
mem[16'h48CC] = 8'h4D;
mem[16'h48CD] = 8'hAD;
mem[16'h48CE] = 8'hB2;
mem[16'h48CF] = 8'h85;
mem[16'h48D0] = 8'hD0;
mem[16'h48D1] = 8'h06;
mem[16'h48D2] = 8'hAD;
mem[16'h48D3] = 8'hB1;
mem[16'h48D4] = 8'h85;
mem[16'h48D5] = 8'h8D;
mem[16'h48D6] = 8'hB0;
mem[16'h48D7] = 8'h85;
mem[16'h48D8] = 8'h60;
mem[16'h48D9] = 8'hA5;
mem[16'h48DA] = 8'h74;
mem[16'h48DB] = 8'hD0;
mem[16'h48DC] = 8'h00;
mem[16'h48DD] = 8'h20;
mem[16'h48DE] = 8'h46;
mem[16'h48DF] = 8'h6D;
mem[16'h48E0] = 8'h20;
mem[16'h48E1] = 8'hCA;
mem[16'h48E2] = 8'h5F;
mem[16'h48E3] = 8'h4C;
mem[16'h48E4] = 8'h0C;
mem[16'h48E5] = 8'h40;
mem[16'h48E6] = 8'h05;
mem[16'h48E7] = 8'hA9;
mem[16'h48E8] = 8'h00;
mem[16'h48E9] = 8'hA0;
mem[16'h48EA] = 8'h80;
mem[16'h48EB] = 8'h20;
mem[16'h48EC] = 8'h86;
mem[16'h48ED] = 8'h68;
mem[16'h48EE] = 8'hA9;
mem[16'h48EF] = 8'h33;
mem[16'h48F0] = 8'h8D;
mem[16'h48F1] = 8'h7F;
mem[16'h48F2] = 8'h68;
mem[16'h48F3] = 8'hAD;
mem[16'h48F4] = 8'hCF;
mem[16'h48F5] = 8'h4D;
mem[16'h48F6] = 8'h85;
mem[16'h48F7] = 8'h57;
mem[16'h48F8] = 8'hAD;
mem[16'h48F9] = 8'hD0;
mem[16'h48FA] = 8'h4D;
mem[16'h48FB] = 8'h85;
mem[16'h48FC] = 8'h56;
mem[16'h48FD] = 8'h20;
mem[16'h48FE] = 8'hE6;
mem[16'h48FF] = 8'h67;
mem[16'h4900] = 8'h60;
mem[16'h4901] = 8'hAE;
mem[16'h4902] = 8'h2E;
mem[16'h4903] = 8'h49;
mem[16'h4904] = 8'hBD;
mem[16'h4905] = 8'h2F;
mem[16'h4906] = 8'h49;
mem[16'h4907] = 8'hBC;
mem[16'h4908] = 8'h34;
mem[16'h4909] = 8'h49;
mem[16'h490A] = 8'h20;
mem[16'h490B] = 8'h86;
mem[16'h490C] = 8'h68;
mem[16'h490D] = 8'hAD;
mem[16'h490E] = 8'hCF;
mem[16'h490F] = 8'h4D;
mem[16'h4910] = 8'h38;
mem[16'h4911] = 8'hE9;
mem[16'h4912] = 8'h03;
mem[16'h4913] = 8'h85;
mem[16'h4914] = 8'h57;
mem[16'h4915] = 8'hAD;
mem[16'h4916] = 8'hD0;
mem[16'h4917] = 8'h4D;
mem[16'h4918] = 8'h38;
mem[16'h4919] = 8'hE9;
mem[16'h491A] = 8'h03;
mem[16'h491B] = 8'h85;
mem[16'h491C] = 8'h56;
mem[16'h491D] = 8'hA9;
mem[16'h491E] = 8'h36;
mem[16'h491F] = 8'h8D;
mem[16'h4920] = 8'h7F;
mem[16'h4921] = 8'h68;
mem[16'h4922] = 8'h20;
mem[16'h4923] = 8'hE6;
mem[16'h4924] = 8'h67;
mem[16'h4925] = 8'hEE;
mem[16'h4926] = 8'h2E;
mem[16'h4927] = 8'h49;
mem[16'h4928] = 8'hA9;
mem[16'h4929] = 8'hFF;
mem[16'h492A] = 8'h20;
mem[16'h492B] = 8'hA8;
mem[16'h492C] = 8'hFC;
mem[16'h492D] = 8'h60;
mem[16'h492E] = 8'hC9;
mem[16'h492F] = 8'h53;
mem[16'h4930] = 8'h89;
mem[16'h4931] = 8'hBF;
mem[16'h4932] = 8'hF5;
mem[16'h4933] = 8'h2B;
mem[16'h4934] = 8'h76;
mem[16'h4935] = 8'h76;
mem[16'h4936] = 8'h76;
mem[16'h4937] = 8'h76;
mem[16'h4938] = 8'h77;
mem[16'h4939] = 8'hA0;
mem[16'h493A] = 8'h64;
mem[16'h493B] = 8'h88;
mem[16'h493C] = 8'hF0;
mem[16'h493D] = 8'h08;
mem[16'h493E] = 8'hA9;
mem[16'h493F] = 8'h64;
mem[16'h4940] = 8'h20;
mem[16'h4941] = 8'hA8;
mem[16'h4942] = 8'hFC;
mem[16'h4943] = 8'h4C;
mem[16'h4944] = 8'h3B;
mem[16'h4945] = 8'h49;
mem[16'h4946] = 8'h60;
mem[16'h4947] = 8'hA0;
mem[16'h4948] = 8'h14;
mem[16'h4949] = 8'h88;
mem[16'h494A] = 8'hF0;
mem[16'h494B] = 8'h08;
mem[16'h494C] = 8'hA9;
mem[16'h494D] = 8'h50;
mem[16'h494E] = 8'h20;
mem[16'h494F] = 8'hA8;
mem[16'h4950] = 8'hFC;
mem[16'h4951] = 8'h4C;
mem[16'h4952] = 8'h49;
mem[16'h4953] = 8'h49;
mem[16'h4954] = 8'h60;
mem[16'h4955] = 8'hA9;
mem[16'h4956] = 8'hC8;
mem[16'h4957] = 8'h8D;
mem[16'h4958] = 8'h22;
mem[16'h4959] = 8'h43;
mem[16'h495A] = 8'hA9;
mem[16'h495B] = 8'h46;
mem[16'h495C] = 8'h8D;
mem[16'h495D] = 8'hB1;
mem[16'h495E] = 8'h85;
mem[16'h495F] = 8'h8D;
mem[16'h4960] = 8'hB0;
mem[16'h4961] = 8'h85;
mem[16'h4962] = 8'hA9;
mem[16'h4963] = 8'h08;
mem[16'h4964] = 8'h8D;
mem[16'h4965] = 8'hAF;
mem[16'h4966] = 8'h4A;
mem[16'h4967] = 8'hA9;
mem[16'h4968] = 8'h03;
mem[16'h4969] = 8'h8D;
mem[16'h496A] = 8'hB1;
mem[16'h496B] = 8'h4A;
mem[16'h496C] = 8'h8D;
mem[16'h496D] = 8'hB3;
mem[16'h496E] = 8'h4A;
mem[16'h496F] = 8'hA9;
mem[16'h4970] = 8'h0E;
mem[16'h4971] = 8'h8D;
mem[16'h4972] = 8'hB0;
mem[16'h4973] = 8'h4A;
mem[16'h4974] = 8'hA9;
mem[16'h4975] = 8'hB4;
mem[16'h4976] = 8'h8D;
mem[16'h4977] = 8'h57;
mem[16'h4978] = 8'h42;
mem[16'h4979] = 8'hA9;
mem[16'h497A] = 8'h64;
mem[16'h497B] = 8'h8D;
mem[16'h497C] = 8'h1F;
mem[16'h497D] = 8'h51;
mem[16'h497E] = 8'hA9;
mem[16'h497F] = 8'h40;
mem[16'h4980] = 8'h8D;
mem[16'h4981] = 8'h0C;
mem[16'h4982] = 8'h54;
mem[16'h4983] = 8'hA9;
mem[16'h4984] = 8'h30;
mem[16'h4985] = 8'h8D;
mem[16'h4986] = 8'h27;
mem[16'h4987] = 8'h53;
mem[16'h4988] = 8'hA9;
mem[16'h4989] = 8'h28;
mem[16'h498A] = 8'h8D;
mem[16'h498B] = 8'hDD;
mem[16'h498C] = 8'h91;
mem[16'h498D] = 8'h8D;
mem[16'h498E] = 8'hDC;
mem[16'h498F] = 8'h91;
mem[16'h4990] = 8'hA9;
mem[16'h4991] = 8'h01;
mem[16'h4992] = 8'h8D;
mem[16'h4993] = 8'hBA;
mem[16'h4994] = 8'h4A;
mem[16'h4995] = 8'h8D;
mem[16'h4996] = 8'hB5;
mem[16'h4997] = 8'h4A;
mem[16'h4998] = 8'h8D;
mem[16'h4999] = 8'hB4;
mem[16'h499A] = 8'h4A;
mem[16'h499B] = 8'h8D;
mem[16'h499C] = 8'hBB;
mem[16'h499D] = 8'h4A;
mem[16'h499E] = 8'h8D;
mem[16'h499F] = 8'hBC;
mem[16'h49A0] = 8'h4A;
mem[16'h49A1] = 8'hA9;
mem[16'h49A2] = 8'h02;
mem[16'h49A3] = 8'h8D;
mem[16'h49A4] = 8'hB2;
mem[16'h49A5] = 8'h4A;
mem[16'h49A6] = 8'h8D;
mem[16'h49A7] = 8'hB8;
mem[16'h49A8] = 8'h4A;
mem[16'h49A9] = 8'h8D;
mem[16'h49AA] = 8'hB9;
mem[16'h49AB] = 8'h4A;
mem[16'h49AC] = 8'h8D;
mem[16'h49AD] = 8'hB6;
mem[16'h49AE] = 8'h4A;
mem[16'h49AF] = 8'h8D;
mem[16'h49B0] = 8'hB7;
mem[16'h49B1] = 8'h4A;
mem[16'h49B2] = 8'h8D;
mem[16'h49B3] = 8'h63;
mem[16'h49B4] = 8'h5E;
mem[16'h49B5] = 8'hA9;
mem[16'h49B6] = 8'h03;
mem[16'h49B7] = 8'h8D;
mem[16'h49B8] = 8'hC4;
mem[16'h49B9] = 8'h5E;
mem[16'h49BA] = 8'hA9;
mem[16'h49BB] = 8'h44;
mem[16'h49BC] = 8'h8D;
mem[16'h49BD] = 8'hAF;
mem[16'h49BE] = 8'h5E;
mem[16'h49BF] = 8'hA9;
mem[16'h49C0] = 8'h28;
mem[16'h49C1] = 8'h8D;
mem[16'h49C2] = 8'h4E;
mem[16'h49C3] = 8'h5E;
mem[16'h49C4] = 8'hA9;
mem[16'h49C5] = 8'h54;
mem[16'h49C6] = 8'h8D;
mem[16'h49C7] = 8'hF8;
mem[16'h49C8] = 8'h5D;
mem[16'h49C9] = 8'hA9;
mem[16'h49CA] = 8'hAA;
mem[16'h49CB] = 8'h8D;
mem[16'h49CC] = 8'hD1;
mem[16'h49CD] = 8'h4F;
mem[16'h49CE] = 8'hA9;
mem[16'h49CF] = 8'hB0;
mem[16'h49D0] = 8'h8D;
mem[16'h49D1] = 8'hE7;
mem[16'h49D2] = 8'h4F;
mem[16'h49D3] = 8'hA9;
mem[16'h49D4] = 8'h4E;
mem[16'h49D5] = 8'h8D;
mem[16'h49D6] = 8'hE3;
mem[16'h49D7] = 8'h51;
mem[16'h49D8] = 8'hA9;
mem[16'h49D9] = 8'hA4;
mem[16'h49DA] = 8'h8D;
mem[16'h49DB] = 8'hF2;
mem[16'h49DC] = 8'h51;
mem[16'h49DD] = 8'hA9;
mem[16'h49DE] = 8'hF4;
mem[16'h49DF] = 8'h8D;
mem[16'h49E0] = 8'h08;
mem[16'h49E1] = 8'h52;
mem[16'h49E2] = 8'hA9;
mem[16'h49E3] = 8'h56;
mem[16'h49E4] = 8'h8D;
mem[16'h49E5] = 8'h6B;
mem[16'h49E6] = 8'h53;
mem[16'h49E7] = 8'hA9;
mem[16'h49E8] = 8'hC0;
mem[16'h49E9] = 8'h8D;
mem[16'h49EA] = 8'h7A;
mem[16'h49EB] = 8'h53;
mem[16'h49EC] = 8'hA9;
mem[16'h49ED] = 8'h62;
mem[16'h49EE] = 8'h8D;
mem[16'h49EF] = 8'hBD;
mem[16'h49F0] = 8'h5F;
mem[16'h49F1] = 8'h8D;
mem[16'h49F2] = 8'hCA;
mem[16'h49F3] = 8'h5D;
mem[16'h49F4] = 8'hA9;
mem[16'h49F5] = 8'h49;
mem[16'h49F6] = 8'h8D;
mem[16'h49F7] = 8'h8F;
mem[16'h49F8] = 8'h5F;
mem[16'h49F9] = 8'h8D;
mem[16'h49FA] = 8'h5E;
mem[16'h49FB] = 8'h5F;
mem[16'h49FC] = 8'hA9;
mem[16'h49FD] = 8'h00;
mem[16'h49FE] = 8'h8D;
mem[16'h49FF] = 8'hC7;
mem[16'h4A00] = 8'h77;
mem[16'h4A01] = 8'h8D;
mem[16'h4A02] = 8'hDF;
mem[16'h4A03] = 8'h91;
mem[16'h4A04] = 8'h8D;
mem[16'h4A05] = 8'hDB;
mem[16'h4A06] = 8'h91;
mem[16'h4A07] = 8'h8D;
mem[16'h4A08] = 8'hDA;
mem[16'h4A09] = 8'h91;
mem[16'h4A0A] = 8'h8D;
mem[16'h4A0B] = 8'hDE;
mem[16'h4A0C] = 8'h91;
mem[16'h4A0D] = 8'h8D;
mem[16'h4A0E] = 8'h5A;
mem[16'h4A0F] = 8'h74;
mem[16'h4A10] = 8'h20;
mem[16'h4A11] = 8'h79;
mem[16'h4A12] = 8'h4A;
mem[16'h4A13] = 8'hA9;
mem[16'h4A14] = 8'h03;
mem[16'h4A15] = 8'h8D;
mem[16'h4A16] = 8'hAA;
mem[16'h4A17] = 8'h4A;
mem[16'h4A18] = 8'h8D;
mem[16'h4A19] = 8'hAB;
mem[16'h4A1A] = 8'h4A;
mem[16'h4A1B] = 8'h8D;
mem[16'h4A1C] = 8'hAC;
mem[16'h4A1D] = 8'h4A;
mem[16'h4A1E] = 8'hA9;
mem[16'h4A1F] = 8'h01;
mem[16'h4A20] = 8'h8D;
mem[16'h4A21] = 8'hAD;
mem[16'h4A22] = 8'h4A;
mem[16'h4A23] = 8'h8D;
mem[16'h4A24] = 8'h23;
mem[16'h4A25] = 8'h43;
mem[16'h4A26] = 8'hA9;
mem[16'h4A27] = 8'h02;
mem[16'h4A28] = 8'h8D;
mem[16'h4A29] = 8'hAE;
mem[16'h4A2A] = 8'h4A;
mem[16'h4A2B] = 8'h8D;
mem[16'h4A2C] = 8'h58;
mem[16'h4A2D] = 8'h42;
mem[16'h4A2E] = 8'hA9;
mem[16'h4A2F] = 8'hD1;
mem[16'h4A30] = 8'h85;
mem[16'h4A31] = 8'h5E;
mem[16'h4A32] = 8'hA9;
mem[16'h4A33] = 8'h4D;
mem[16'h4A34] = 8'h85;
mem[16'h4A35] = 8'h5F;
mem[16'h4A36] = 8'hAD;
mem[16'h4A37] = 8'hCE;
mem[16'h4A38] = 8'h44;
mem[16'h4A39] = 8'hC9;
mem[16'h4A3A] = 8'h01;
mem[16'h4A3B] = 8'hF0;
mem[16'h4A3C] = 8'h39;
mem[16'h4A3D] = 8'hA9;
mem[16'h4A3E] = 8'h03;
mem[16'h4A3F] = 8'h8D;
mem[16'h4A40] = 8'hCD;
mem[16'h4A41] = 8'h6A;
mem[16'h4A42] = 8'h8D;
mem[16'h4A43] = 8'h88;
mem[16'h4A44] = 8'h6B;
mem[16'h4A45] = 8'hA9;
mem[16'h4A46] = 8'h33;
mem[16'h4A47] = 8'h8D;
mem[16'h4A48] = 8'hC9;
mem[16'h4A49] = 8'h77;
mem[16'h4A4A] = 8'h8D;
mem[16'h4A4B] = 8'hCB;
mem[16'h4A4C] = 8'h77;
mem[16'h4A4D] = 8'hA9;
mem[16'h4A4E] = 8'h02;
mem[16'h4A4F] = 8'h8D;
mem[16'h4A50] = 8'hB1;
mem[16'h4A51] = 8'h4A;
mem[16'h4A52] = 8'h8D;
mem[16'h4A53] = 8'hC7;
mem[16'h4A54] = 8'h77;
mem[16'h4A55] = 8'hA9;
mem[16'h4A56] = 8'h01;
mem[16'h4A57] = 8'h8D;
mem[16'h4A58] = 8'h5A;
mem[16'h4A59] = 8'h74;
mem[16'h4A5A] = 8'hA9;
mem[16'h4A5B] = 8'h0A;
mem[16'h4A5C] = 8'h8D;
mem[16'h4A5D] = 8'hDF;
mem[16'h4A5E] = 8'h91;
mem[16'h4A5F] = 8'h8D;
mem[16'h4A60] = 8'hDE;
mem[16'h4A61] = 8'h91;
mem[16'h4A62] = 8'hA9;
mem[16'h4A63] = 8'h01;
mem[16'h4A64] = 8'h8D;
mem[16'h4A65] = 8'hB2;
mem[16'h4A66] = 8'h4A;
mem[16'h4A67] = 8'hA9;
mem[16'h4A68] = 8'h78;
mem[16'h4A69] = 8'h8D;
mem[16'h4A6A] = 8'h6B;
mem[16'h4A6B] = 8'h53;
mem[16'h4A6C] = 8'hA9;
mem[16'h4A6D] = 8'hA0;
mem[16'h4A6E] = 8'h8D;
mem[16'h4A6F] = 8'h1F;
mem[16'h4A70] = 8'h51;
mem[16'h4A71] = 8'hA9;
mem[16'h4A72] = 8'hC8;
mem[16'h4A73] = 8'h8D;
mem[16'h4A74] = 8'hD1;
mem[16'h4A75] = 8'h4F;
mem[16'h4A76] = 8'h4C;
mem[16'h4A77] = 8'h18;
mem[16'h4A78] = 8'h40;
mem[16'h4A79] = 8'hA9;
mem[16'h4A7A] = 8'h00;
mem[16'h4A7B] = 8'h8D;
mem[16'h4A7C] = 8'hD9;
mem[16'h4A7D] = 8'h77;
mem[16'h4A7E] = 8'h85;
mem[16'h4A7F] = 8'h8B;
mem[16'h4A80] = 8'h8D;
mem[16'h4A81] = 8'hB2;
mem[16'h4A82] = 8'h85;
mem[16'h4A83] = 8'h8D;
mem[16'h4A84] = 8'h33;
mem[16'h4A85] = 8'h7B;
mem[16'h4A86] = 8'h8D;
mem[16'h4A87] = 8'hC2;
mem[16'h4A88] = 8'h62;
mem[16'h4A89] = 8'h8D;
mem[16'h4A8A] = 8'hC1;
mem[16'h4A8B] = 8'h62;
mem[16'h4A8C] = 8'h8D;
mem[16'h4A8D] = 8'hC3;
mem[16'h4A8E] = 8'h62;
mem[16'h4A8F] = 8'h8D;
mem[16'h4A90] = 8'hC0;
mem[16'h4A91] = 8'h62;
mem[16'h4A92] = 8'h8D;
mem[16'h4A93] = 8'hD8;
mem[16'h4A94] = 8'h77;
mem[16'h4A95] = 8'h85;
mem[16'h4A96] = 8'h87;
mem[16'h4A97] = 8'hA2;
mem[16'h4A98] = 8'h0E;
mem[16'h4A99] = 8'hCA;
mem[16'h4A9A] = 8'h30;
mem[16'h4A9B] = 8'h0D;
mem[16'h4A9C] = 8'hA9;
mem[16'h4A9D] = 8'h00;
mem[16'h4A9E] = 8'h9D;
mem[16'h4A9F] = 8'h75;
mem[16'h4AA0] = 8'h5B;
mem[16'h4AA1] = 8'hA9;
mem[16'h4AA2] = 8'h07;
mem[16'h4AA3] = 8'h9D;
mem[16'h4AA4] = 8'h83;
mem[16'h4AA5] = 8'h5B;
mem[16'h4AA6] = 8'h4C;
mem[16'h4AA7] = 8'h99;
mem[16'h4AA8] = 8'h4A;
mem[16'h4AA9] = 8'h60;
mem[16'h4AAA] = 8'h03;
mem[16'h4AAB] = 8'h03;
mem[16'h4AAC] = 8'h03;
mem[16'h4AAD] = 8'h01;
mem[16'h4AAE] = 8'h02;
mem[16'h4AAF] = 8'h08;
mem[16'h4AB0] = 8'h0E;
mem[16'h4AB1] = 8'h03;
mem[16'h4AB2] = 8'h02;
mem[16'h4AB3] = 8'h03;
mem[16'h4AB4] = 8'h01;
mem[16'h4AB5] = 8'h01;
mem[16'h4AB6] = 8'h02;
mem[16'h4AB7] = 8'h02;
mem[16'h4AB8] = 8'h02;
mem[16'h4AB9] = 8'h02;
mem[16'h4ABA] = 8'h01;
mem[16'h4ABB] = 8'h01;
mem[16'h4ABC] = 8'h01;
mem[16'h4ABD] = 8'hA5;
mem[16'h4ABE] = 8'h87;
mem[16'h4ABF] = 8'hF0;
mem[16'h4AC0] = 8'h03;
mem[16'h4AC1] = 8'h4C;
mem[16'h4AC2] = 8'h55;
mem[16'h4AC3] = 8'h4B;
mem[16'h4AC4] = 8'hA5;
mem[16'h4AC5] = 8'h85;
mem[16'h4AC6] = 8'hF0;
mem[16'h4AC7] = 8'h03;
mem[16'h4AC8] = 8'h20;
mem[16'h4AC9] = 8'h52;
mem[16'h4ACA] = 8'h7F;
mem[16'h4ACB] = 8'hAD;
mem[16'h4ACC] = 8'h00;
mem[16'h4ACD] = 8'hC0;
mem[16'h4ACE] = 8'hC5;
mem[16'h4ACF] = 8'h7D;
mem[16'h4AD0] = 8'hD0;
mem[16'h4AD1] = 8'h1C;
mem[16'h4AD2] = 8'h85;
mem[16'h4AD3] = 8'h88;
mem[16'h4AD4] = 8'hAD;
mem[16'h4AD5] = 8'h10;
mem[16'h4AD6] = 8'hC0;
mem[16'h4AD7] = 8'hA9;
mem[16'h4AD8] = 8'h01;
mem[16'h4AD9] = 8'h85;
mem[16'h4ADA] = 8'h87;
mem[16'h4ADB] = 8'h20;
mem[16'h4ADC] = 8'hD9;
mem[16'h4ADD] = 8'h4C;
mem[16'h4ADE] = 8'hAD;
mem[16'h4ADF] = 8'hD0;
mem[16'h4AE0] = 8'h4D;
mem[16'h4AE1] = 8'h38;
mem[16'h4AE2] = 8'hE9;
mem[16'h4AE3] = 8'h07;
mem[16'h4AE4] = 8'h8D;
mem[16'h4AE5] = 8'hD0;
mem[16'h4AE6] = 8'h4D;
mem[16'h4AE7] = 8'h20;
mem[16'h4AE8] = 8'h0D;
mem[16'h4AE9] = 8'h4D;
mem[16'h4AEA] = 8'h20;
mem[16'h4AEB] = 8'h95;
mem[16'h4AEC] = 8'h4C;
mem[16'h4AED] = 8'h60;
mem[16'h4AEE] = 8'hC5;
mem[16'h4AEF] = 8'h7E;
mem[16'h4AF0] = 8'hD0;
mem[16'h4AF1] = 8'h23;
mem[16'h4AF2] = 8'h85;
mem[16'h4AF3] = 8'h88;
mem[16'h4AF4] = 8'hAD;
mem[16'h4AF5] = 8'h10;
mem[16'h4AF6] = 8'hC0;
mem[16'h4AF7] = 8'hAD;
mem[16'h4AF8] = 8'hD0;
mem[16'h4AF9] = 8'h4D;
mem[16'h4AFA] = 8'hC9;
mem[16'h4AFB] = 8'hAF;
mem[16'h4AFC] = 8'hF0;
mem[16'h4AFD] = 8'h56;
mem[16'h4AFE] = 8'hA9;
mem[16'h4AFF] = 8'h01;
mem[16'h4B00] = 8'h85;
mem[16'h4B01] = 8'h87;
mem[16'h4B02] = 8'h20;
mem[16'h4B03] = 8'hD9;
mem[16'h4B04] = 8'h4C;
mem[16'h4B05] = 8'hAD;
mem[16'h4B06] = 8'hD0;
mem[16'h4B07] = 8'h4D;
mem[16'h4B08] = 8'h18;
mem[16'h4B09] = 8'h69;
mem[16'h4B0A] = 8'h07;
mem[16'h4B0B] = 8'h8D;
mem[16'h4B0C] = 8'hD0;
mem[16'h4B0D] = 8'h4D;
mem[16'h4B0E] = 8'h20;
mem[16'h4B0F] = 8'h45;
mem[16'h4B10] = 8'h4D;
mem[16'h4B11] = 8'h20;
mem[16'h4B12] = 8'h95;
mem[16'h4B13] = 8'h4C;
mem[16'h4B14] = 8'h60;
mem[16'h4B15] = 8'hC5;
mem[16'h4B16] = 8'h7F;
mem[16'h4B17] = 8'hD0;
mem[16'h4B18] = 8'h1C;
mem[16'h4B19] = 8'h85;
mem[16'h4B1A] = 8'h88;
mem[16'h4B1B] = 8'hAD;
mem[16'h4B1C] = 8'h10;
mem[16'h4B1D] = 8'hC0;
mem[16'h4B1E] = 8'hA9;
mem[16'h4B1F] = 8'h01;
mem[16'h4B20] = 8'h85;
mem[16'h4B21] = 8'h87;
mem[16'h4B22] = 8'h20;
mem[16'h4B23] = 8'hD9;
mem[16'h4B24] = 8'h4C;
mem[16'h4B25] = 8'hAD;
mem[16'h4B26] = 8'hCF;
mem[16'h4B27] = 8'h4D;
mem[16'h4B28] = 8'h38;
mem[16'h4B29] = 8'hE9;
mem[16'h4B2A] = 8'h05;
mem[16'h4B2B] = 8'h8D;
mem[16'h4B2C] = 8'hCF;
mem[16'h4B2D] = 8'h4D;
mem[16'h4B2E] = 8'h20;
mem[16'h4B2F] = 8'h27;
mem[16'h4B30] = 8'h4D;
mem[16'h4B31] = 8'h20;
mem[16'h4B32] = 8'h95;
mem[16'h4B33] = 8'h4C;
mem[16'h4B34] = 8'h60;
mem[16'h4B35] = 8'hC5;
mem[16'h4B36] = 8'h80;
mem[16'h4B37] = 8'hD0;
mem[16'h4B38] = 8'h1B;
mem[16'h4B39] = 8'h85;
mem[16'h4B3A] = 8'h88;
mem[16'h4B3B] = 8'hAD;
mem[16'h4B3C] = 8'h10;
mem[16'h4B3D] = 8'hC0;
mem[16'h4B3E] = 8'hA9;
mem[16'h4B3F] = 8'h01;
mem[16'h4B40] = 8'h85;
mem[16'h4B41] = 8'h87;
mem[16'h4B42] = 8'h20;
mem[16'h4B43] = 8'hD9;
mem[16'h4B44] = 8'h4C;
mem[16'h4B45] = 8'hAD;
mem[16'h4B46] = 8'hCF;
mem[16'h4B47] = 8'h4D;
mem[16'h4B48] = 8'h18;
mem[16'h4B49] = 8'h69;
mem[16'h4B4A] = 8'h05;
mem[16'h4B4B] = 8'h8D;
mem[16'h4B4C] = 8'hCF;
mem[16'h4B4D] = 8'h4D;
mem[16'h4B4E] = 8'h20;
mem[16'h4B4F] = 8'h36;
mem[16'h4B50] = 8'h4D;
mem[16'h4B51] = 8'h20;
mem[16'h4B52] = 8'h95;
mem[16'h4B53] = 8'h4C;
mem[16'h4B54] = 8'h60;
mem[16'h4B55] = 8'hAD;
mem[16'h4B56] = 8'h10;
mem[16'h4B57] = 8'hC0;
mem[16'h4B58] = 8'hA5;
mem[16'h4B59] = 8'h88;
mem[16'h4B5A] = 8'hC5;
mem[16'h4B5B] = 8'h7D;
mem[16'h4B5C] = 8'hD0;
mem[16'h4B5D] = 8'h25;
mem[16'h4B5E] = 8'h20;
mem[16'h4B5F] = 8'h0D;
mem[16'h4B60] = 8'h4D;
mem[16'h4B61] = 8'hAD;
mem[16'h4B62] = 8'hD0;
mem[16'h4B63] = 8'h4D;
mem[16'h4B64] = 8'h38;
mem[16'h4B65] = 8'hE9;
mem[16'h4B66] = 8'h07;
mem[16'h4B67] = 8'h8D;
mem[16'h4B68] = 8'hD0;
mem[16'h4B69] = 8'h4D;
mem[16'h4B6A] = 8'hC6;
mem[16'h4B6B] = 8'h87;
mem[16'h4B6C] = 8'h20;
mem[16'h4B6D] = 8'h95;
mem[16'h4B6E] = 8'h4C;
mem[16'h4B6F] = 8'hA5;
mem[16'h4B70] = 8'h87;
mem[16'h4B71] = 8'hF0;
mem[16'h4B72] = 8'h04;
mem[16'h4B73] = 8'h20;
mem[16'h4B74] = 8'h0D;
mem[16'h4B75] = 8'h4D;
mem[16'h4B76] = 8'h60;
mem[16'h4B77] = 8'h20;
mem[16'h4B78] = 8'hD9;
mem[16'h4B79] = 8'h4C;
mem[16'h4B7A] = 8'hA9;
mem[16'h4B7B] = 8'h10;
mem[16'h4B7C] = 8'h20;
mem[16'h4B7D] = 8'h89;
mem[16'h4B7E] = 8'h66;
mem[16'h4B7F] = 8'h20;
mem[16'h4B80] = 8'h59;
mem[16'h4B81] = 8'h43;
mem[16'h4B82] = 8'h60;
mem[16'h4B83] = 8'hC5;
mem[16'h4B84] = 8'h7E;
mem[16'h4B85] = 8'hD0;
mem[16'h4B86] = 8'h20;
mem[16'h4B87] = 8'h20;
mem[16'h4B88] = 8'h45;
mem[16'h4B89] = 8'h4D;
mem[16'h4B8A] = 8'hAD;
mem[16'h4B8B] = 8'hD0;
mem[16'h4B8C] = 8'h4D;
mem[16'h4B8D] = 8'h18;
mem[16'h4B8E] = 8'h69;
mem[16'h4B8F] = 8'h07;
mem[16'h4B90] = 8'h8D;
mem[16'h4B91] = 8'hD0;
mem[16'h4B92] = 8'h4D;
mem[16'h4B93] = 8'hC6;
mem[16'h4B94] = 8'h87;
mem[16'h4B95] = 8'h20;
mem[16'h4B96] = 8'h95;
mem[16'h4B97] = 8'h4C;
mem[16'h4B98] = 8'hA5;
mem[16'h4B99] = 8'h87;
mem[16'h4B9A] = 8'hF0;
mem[16'h4B9B] = 8'h04;
mem[16'h4B9C] = 8'h20;
mem[16'h4B9D] = 8'h45;
mem[16'h4B9E] = 8'h4D;
mem[16'h4B9F] = 8'h60;
mem[16'h4BA0] = 8'h20;
mem[16'h4BA1] = 8'hD9;
mem[16'h4BA2] = 8'h4C;
mem[16'h4BA3] = 8'h20;
mem[16'h4BA4] = 8'h59;
mem[16'h4BA5] = 8'h43;
mem[16'h4BA6] = 8'h60;
mem[16'h4BA7] = 8'hC5;
mem[16'h4BA8] = 8'h7F;
mem[16'h4BA9] = 8'hD0;
mem[16'h4BAA] = 8'h20;
mem[16'h4BAB] = 8'h20;
mem[16'h4BAC] = 8'h27;
mem[16'h4BAD] = 8'h4D;
mem[16'h4BAE] = 8'hAD;
mem[16'h4BAF] = 8'hCF;
mem[16'h4BB0] = 8'h4D;
mem[16'h4BB1] = 8'h38;
mem[16'h4BB2] = 8'hE9;
mem[16'h4BB3] = 8'h05;
mem[16'h4BB4] = 8'h8D;
mem[16'h4BB5] = 8'hCF;
mem[16'h4BB6] = 8'h4D;
mem[16'h4BB7] = 8'hC6;
mem[16'h4BB8] = 8'h87;
mem[16'h4BB9] = 8'h20;
mem[16'h4BBA] = 8'h95;
mem[16'h4BBB] = 8'h4C;
mem[16'h4BBC] = 8'hA5;
mem[16'h4BBD] = 8'h87;
mem[16'h4BBE] = 8'hF0;
mem[16'h4BBF] = 8'h04;
mem[16'h4BC0] = 8'h20;
mem[16'h4BC1] = 8'h27;
mem[16'h4BC2] = 8'h4D;
mem[16'h4BC3] = 8'h60;
mem[16'h4BC4] = 8'h20;
mem[16'h4BC5] = 8'hD9;
mem[16'h4BC6] = 8'h4C;
mem[16'h4BC7] = 8'h20;
mem[16'h4BC8] = 8'h59;
mem[16'h4BC9] = 8'h43;
mem[16'h4BCA] = 8'h60;
mem[16'h4BCB] = 8'hC5;
mem[16'h4BCC] = 8'h80;
mem[16'h4BCD] = 8'hD0;
mem[16'h4BCE] = 8'h1F;
mem[16'h4BCF] = 8'h20;
mem[16'h4BD0] = 8'h36;
mem[16'h4BD1] = 8'h4D;
mem[16'h4BD2] = 8'hAD;
mem[16'h4BD3] = 8'hCF;
mem[16'h4BD4] = 8'h4D;
mem[16'h4BD5] = 8'h18;
mem[16'h4BD6] = 8'h69;
mem[16'h4BD7] = 8'h05;
mem[16'h4BD8] = 8'h8D;
mem[16'h4BD9] = 8'hCF;
mem[16'h4BDA] = 8'h4D;
mem[16'h4BDB] = 8'hC6;
mem[16'h4BDC] = 8'h87;
mem[16'h4BDD] = 8'h20;
mem[16'h4BDE] = 8'h95;
mem[16'h4BDF] = 8'h4C;
mem[16'h4BE0] = 8'hA5;
mem[16'h4BE1] = 8'h87;
mem[16'h4BE2] = 8'hF0;
mem[16'h4BE3] = 8'h04;
mem[16'h4BE4] = 8'h20;
mem[16'h4BE5] = 8'h36;
mem[16'h4BE6] = 8'h4D;
mem[16'h4BE7] = 8'h60;
mem[16'h4BE8] = 8'h20;
mem[16'h4BE9] = 8'hD9;
mem[16'h4BEA] = 8'h4C;
mem[16'h4BEB] = 8'h20;
mem[16'h4BEC] = 8'h59;
mem[16'h4BED] = 8'h43;
mem[16'h4BEE] = 8'h60;
mem[16'h4BEF] = 8'hA9;
mem[16'h4BF0] = 8'hFD;
mem[16'h4BF1] = 8'h85;
mem[16'h4BF2] = 8'h55;
mem[16'h4BF3] = 8'hA9;
mem[16'h4BF4] = 8'h50;
mem[16'h4BF5] = 8'h85;
mem[16'h4BF6] = 8'h50;
mem[16'h4BF7] = 8'hA9;
mem[16'h4BF8] = 8'h04;
mem[16'h4BF9] = 8'h85;
mem[16'h4BFA] = 8'h52;
mem[16'h4BFB] = 8'h85;
mem[16'h4BFC] = 8'h53;
mem[16'h4BFD] = 8'h20;
mem[16'h4BFE] = 8'h00;
mem[16'h4BFF] = 8'h65;
mem[16'h4C00] = 8'hA5;
mem[16'h4C01] = 8'h50;
mem[16'h4C02] = 8'h38;
mem[16'h4C03] = 8'hE9;
mem[16'h4C04] = 8'h14;
mem[16'h4C05] = 8'h85;
mem[16'h4C06] = 8'h50;
mem[16'h4C07] = 8'hC9;
mem[16'h4C08] = 8'h14;
mem[16'h4C09] = 8'hD0;
mem[16'h4C0A] = 8'hEC;
mem[16'h4C0B] = 8'h60;
mem[16'h4C0C] = 8'hA9;
mem[16'h4C0D] = 8'h00;
mem[16'h4C0E] = 8'h85;
mem[16'h4C0F] = 8'h55;
mem[16'h4C10] = 8'hAD;
mem[16'h4C11] = 8'h22;
mem[16'h4C12] = 8'h4C;
mem[16'h4C13] = 8'h85;
mem[16'h4C14] = 8'h50;
mem[16'h4C15] = 8'hA9;
mem[16'h4C16] = 8'h08;
mem[16'h4C17] = 8'h85;
mem[16'h4C18] = 8'h52;
mem[16'h4C19] = 8'h85;
mem[16'h4C1A] = 8'h53;
mem[16'h4C1B] = 8'h20;
mem[16'h4C1C] = 8'h00;
mem[16'h4C1D] = 8'h65;
mem[16'h4C1E] = 8'hCE;
mem[16'h4C1F] = 8'h22;
mem[16'h4C20] = 8'h4C;
mem[16'h4C21] = 8'h60;
mem[16'h4C22] = 8'h00;
mem[16'h4C23] = 8'hA9;
mem[16'h4C24] = 8'h00;
mem[16'h4C25] = 8'h85;
mem[16'h4C26] = 8'h55;
mem[16'h4C27] = 8'hA9;
mem[16'h4C28] = 8'h14;
mem[16'h4C29] = 8'h8D;
mem[16'h4C2A] = 8'h6C;
mem[16'h4C2B] = 8'h4C;
mem[16'h4C2C] = 8'hA9;
mem[16'h4C2D] = 8'h12;
mem[16'h4C2E] = 8'h85;
mem[16'h4C2F] = 8'h50;
mem[16'h4C30] = 8'hA9;
mem[16'h4C31] = 8'h0C;
mem[16'h4C32] = 8'h85;
mem[16'h4C33] = 8'h52;
mem[16'h4C34] = 8'h85;
mem[16'h4C35] = 8'h53;
mem[16'h4C36] = 8'h20;
mem[16'h4C37] = 8'h00;
mem[16'h4C38] = 8'h65;
mem[16'h4C39] = 8'hA5;
mem[16'h4C3A] = 8'h50;
mem[16'h4C3B] = 8'h49;
mem[16'h4C3C] = 8'h06;
mem[16'h4C3D] = 8'h85;
mem[16'h4C3E] = 8'h50;
mem[16'h4C3F] = 8'hA9;
mem[16'h4C40] = 8'h64;
mem[16'h4C41] = 8'h20;
mem[16'h4C42] = 8'hA8;
mem[16'h4C43] = 8'hFC;
mem[16'h4C44] = 8'hCE;
mem[16'h4C45] = 8'h6C;
mem[16'h4C46] = 8'h4C;
mem[16'h4C47] = 8'hD0;
mem[16'h4C48] = 8'hE7;
mem[16'h4C49] = 8'h60;
mem[16'h4C4A] = 8'hA9;
mem[16'h4C4B] = 8'hFD;
mem[16'h4C4C] = 8'h85;
mem[16'h4C4D] = 8'h55;
mem[16'h4C4E] = 8'hA9;
mem[16'h4C4F] = 8'h04;
mem[16'h4C50] = 8'h8D;
mem[16'h4C51] = 8'h6C;
mem[16'h4C52] = 8'h4C;
mem[16'h4C53] = 8'hA9;
mem[16'h4C54] = 8'h10;
mem[16'h4C55] = 8'h85;
mem[16'h4C56] = 8'h50;
mem[16'h4C57] = 8'hA9;
mem[16'h4C58] = 8'h04;
mem[16'h4C59] = 8'h85;
mem[16'h4C5A] = 8'h52;
mem[16'h4C5B] = 8'h85;
mem[16'h4C5C] = 8'h53;
mem[16'h4C5D] = 8'h20;
mem[16'h4C5E] = 8'h00;
mem[16'h4C5F] = 8'h65;
mem[16'h4C60] = 8'hA5;
mem[16'h4C61] = 8'h50;
mem[16'h4C62] = 8'h49;
mem[16'h4C63] = 8'h20;
mem[16'h4C64] = 8'h85;
mem[16'h4C65] = 8'h50;
mem[16'h4C66] = 8'hCE;
mem[16'h4C67] = 8'h6C;
mem[16'h4C68] = 8'h4C;
mem[16'h4C69] = 8'hD0;
mem[16'h4C6A] = 8'hEC;
mem[16'h4C6B] = 8'h60;
mem[16'h4C6C] = 8'h00;
mem[16'h4C6D] = 8'hA9;
mem[16'h4C6E] = 8'h00;
mem[16'h4C6F] = 8'h85;
mem[16'h4C70] = 8'h55;
mem[16'h4C71] = 8'hA9;
mem[16'h4C72] = 8'h14;
mem[16'h4C73] = 8'h8D;
mem[16'h4C74] = 8'h6C;
mem[16'h4C75] = 8'h4C;
mem[16'h4C76] = 8'hA9;
mem[16'h4C77] = 8'hA0;
mem[16'h4C78] = 8'h85;
mem[16'h4C79] = 8'h50;
mem[16'h4C7A] = 8'hA9;
mem[16'h4C7B] = 8'h0C;
mem[16'h4C7C] = 8'h85;
mem[16'h4C7D] = 8'h52;
mem[16'h4C7E] = 8'h85;
mem[16'h4C7F] = 8'h53;
mem[16'h4C80] = 8'h20;
mem[16'h4C81] = 8'h00;
mem[16'h4C82] = 8'h65;
mem[16'h4C83] = 8'hA5;
mem[16'h4C84] = 8'h50;
mem[16'h4C85] = 8'h49;
mem[16'h4C86] = 8'h20;
mem[16'h4C87] = 8'h85;
mem[16'h4C88] = 8'h50;
mem[16'h4C89] = 8'hA9;
mem[16'h4C8A] = 8'h50;
mem[16'h4C8B] = 8'h20;
mem[16'h4C8C] = 8'hA8;
mem[16'h4C8D] = 8'hFC;
mem[16'h4C8E] = 8'hCE;
mem[16'h4C8F] = 8'h6C;
mem[16'h4C90] = 8'h4C;
mem[16'h4C91] = 8'hD0;
mem[16'h4C92] = 8'hE7;
mem[16'h4C93] = 8'h60;
mem[16'h4C94] = 8'h00;
mem[16'h4C95] = 8'hA6;
mem[16'h4C96] = 8'h87;
mem[16'h4C97] = 8'hBD;
mem[16'h4C98] = 8'hAA;
mem[16'h4C99] = 8'h4C;
mem[16'h4C9A] = 8'h85;
mem[16'h4C9B] = 8'h50;
mem[16'h4C9C] = 8'hA9;
mem[16'h4C9D] = 8'h00;
mem[16'h4C9E] = 8'h85;
mem[16'h4C9F] = 8'h55;
mem[16'h4CA0] = 8'hA9;
mem[16'h4CA1] = 8'h02;
mem[16'h4CA2] = 8'h85;
mem[16'h4CA3] = 8'h52;
mem[16'h4CA4] = 8'h85;
mem[16'h4CA5] = 8'h53;
mem[16'h4CA6] = 8'h20;
mem[16'h4CA7] = 8'h00;
mem[16'h4CA8] = 8'h65;
mem[16'h4CA9] = 8'h60;
mem[16'h4CAA] = 8'h16;
mem[16'h4CAB] = 8'h11;
mem[16'h4CAC] = 8'h10;
mem[16'h4CAD] = 8'h11;
mem[16'h4CAE] = 8'hA5;
mem[16'h4CAF] = 8'h87;
mem[16'h4CB0] = 8'hD0;
mem[16'h4CB1] = 8'h04;
mem[16'h4CB2] = 8'h20;
mem[16'h4CB3] = 8'hD9;
mem[16'h4CB4] = 8'h4C;
mem[16'h4CB5] = 8'h60;
mem[16'h4CB6] = 8'hA5;
mem[16'h4CB7] = 8'h88;
mem[16'h4CB8] = 8'hC5;
mem[16'h4CB9] = 8'h7D;
mem[16'h4CBA] = 8'hD0;
mem[16'h4CBB] = 8'h04;
mem[16'h4CBC] = 8'h20;
mem[16'h4CBD] = 8'h0D;
mem[16'h4CBE] = 8'h4D;
mem[16'h4CBF] = 8'h60;
mem[16'h4CC0] = 8'hC5;
mem[16'h4CC1] = 8'h7E;
mem[16'h4CC2] = 8'hD0;
mem[16'h4CC3] = 8'h04;
mem[16'h4CC4] = 8'h20;
mem[16'h4CC5] = 8'h45;
mem[16'h4CC6] = 8'h4D;
mem[16'h4CC7] = 8'h60;
mem[16'h4CC8] = 8'hC5;
mem[16'h4CC9] = 8'h7F;
mem[16'h4CCA] = 8'hD0;
mem[16'h4CCB] = 8'h04;
mem[16'h4CCC] = 8'h20;
mem[16'h4CCD] = 8'h27;
mem[16'h4CCE] = 8'h4D;
mem[16'h4CCF] = 8'h60;
mem[16'h4CD0] = 8'hC5;
mem[16'h4CD1] = 8'h80;
mem[16'h4CD2] = 8'hD0;
mem[16'h4CD3] = 8'h03;
mem[16'h4CD4] = 8'h20;
mem[16'h4CD5] = 8'h36;
mem[16'h4CD6] = 8'h4D;
mem[16'h4CD7] = 8'h60;
mem[16'h4CD8] = 8'h60;
mem[16'h4CD9] = 8'hAD;
mem[16'h4CDA] = 8'hD0;
mem[16'h4CDB] = 8'h4D;
mem[16'h4CDC] = 8'h85;
mem[16'h4CDD] = 8'h56;
mem[16'h4CDE] = 8'hA9;
mem[16'h4CDF] = 8'hF3;
mem[16'h4CE0] = 8'hA0;
mem[16'h4CE1] = 8'h4C;
mem[16'h4CE2] = 8'h20;
mem[16'h4CE3] = 8'h42;
mem[16'h4CE4] = 8'h6A;
mem[16'h4CE5] = 8'hA9;
mem[16'h4CE6] = 8'h1A;
mem[16'h4CE7] = 8'h8D;
mem[16'h4CE8] = 8'hF9;
mem[16'h4CE9] = 8'h69;
mem[16'h4CEA] = 8'hAD;
mem[16'h4CEB] = 8'hCF;
mem[16'h4CEC] = 8'h4D;
mem[16'h4CED] = 8'h85;
mem[16'h4CEE] = 8'h57;
mem[16'h4CEF] = 8'h20;
mem[16'h4CF0] = 8'h33;
mem[16'h4CF1] = 8'h69;
mem[16'h4CF2] = 8'h60;
mem[16'h4CF3] = 8'h00;
mem[16'h4CF4] = 8'h00;
mem[16'h4CF5] = 8'h40;
mem[16'h4CF6] = 8'h01;
mem[16'h4CF7] = 8'h60;
mem[16'h4CF8] = 8'h03;
mem[16'h4CF9] = 8'h60;
mem[16'h4CFA] = 8'h03;
mem[16'h4CFB] = 8'h40;
mem[16'h4CFC] = 8'h01;
mem[16'h4CFD] = 8'h60;
mem[16'h4CFE] = 8'h03;
mem[16'h4CFF] = 8'h70;
mem[16'h4D00] = 8'h07;
mem[16'h4D01] = 8'h74;
mem[16'h4D02] = 8'h17;
mem[16'h4D03] = 8'h7C;
mem[16'h4D04] = 8'h1F;
mem[16'h4D05] = 8'h7C;
mem[16'h4D06] = 8'h1F;
mem[16'h4D07] = 8'h44;
mem[16'h4D08] = 8'h12;
mem[16'h4D09] = 8'h0E;
mem[16'h4D0A] = 8'h38;
mem[16'h4D0B] = 8'h0E;
mem[16'h4D0C] = 8'h38;
mem[16'h4D0D] = 8'hA9;
mem[16'h4D0E] = 8'h54;
mem[16'h4D0F] = 8'hA0;
mem[16'h4D10] = 8'h4D;
mem[16'h4D11] = 8'h20;
mem[16'h4D12] = 8'h42;
mem[16'h4D13] = 8'h6A;
mem[16'h4D14] = 8'hA9;
mem[16'h4D15] = 8'h1A;
mem[16'h4D16] = 8'h8D;
mem[16'h4D17] = 8'hF9;
mem[16'h4D18] = 8'h69;
mem[16'h4D19] = 8'hAD;
mem[16'h4D1A] = 8'hCF;
mem[16'h4D1B] = 8'h4D;
mem[16'h4D1C] = 8'h85;
mem[16'h4D1D] = 8'h57;
mem[16'h4D1E] = 8'hAD;
mem[16'h4D1F] = 8'hD0;
mem[16'h4D20] = 8'h4D;
mem[16'h4D21] = 8'h85;
mem[16'h4D22] = 8'h56;
mem[16'h4D23] = 8'h20;
mem[16'h4D24] = 8'h33;
mem[16'h4D25] = 8'h69;
mem[16'h4D26] = 8'h60;
mem[16'h4D27] = 8'hA9;
mem[16'h4D28] = 8'h88;
mem[16'h4D29] = 8'hA0;
mem[16'h4D2A] = 8'h4D;
mem[16'h4D2B] = 8'h20;
mem[16'h4D2C] = 8'h42;
mem[16'h4D2D] = 8'h6A;
mem[16'h4D2E] = 8'hA9;
mem[16'h4D2F] = 8'h16;
mem[16'h4D30] = 8'h8D;
mem[16'h4D31] = 8'hF9;
mem[16'h4D32] = 8'h69;
mem[16'h4D33] = 8'h4C;
mem[16'h4D34] = 8'h19;
mem[16'h4D35] = 8'h4D;
mem[16'h4D36] = 8'hA9;
mem[16'h4D37] = 8'h9E;
mem[16'h4D38] = 8'hA0;
mem[16'h4D39] = 8'h4D;
mem[16'h4D3A] = 8'h20;
mem[16'h4D3B] = 8'h42;
mem[16'h4D3C] = 8'h6A;
mem[16'h4D3D] = 8'hA9;
mem[16'h4D3E] = 8'h16;
mem[16'h4D3F] = 8'h8D;
mem[16'h4D40] = 8'hF9;
mem[16'h4D41] = 8'h69;
mem[16'h4D42] = 8'h4C;
mem[16'h4D43] = 8'h19;
mem[16'h4D44] = 8'h4D;
mem[16'h4D45] = 8'hA9;
mem[16'h4D46] = 8'h6E;
mem[16'h4D47] = 8'hA0;
mem[16'h4D48] = 8'h4D;
mem[16'h4D49] = 8'h20;
mem[16'h4D4A] = 8'h42;
mem[16'h4D4B] = 8'h6A;
mem[16'h4D4C] = 8'hA9;
mem[16'h4D4D] = 8'h1A;
mem[16'h4D4E] = 8'h8D;
mem[16'h4D4F] = 8'hF9;
mem[16'h4D50] = 8'h69;
mem[16'h4D51] = 8'h4C;
mem[16'h4D52] = 8'h19;
mem[16'h4D53] = 8'h4D;
mem[16'h4D54] = 8'h60;
mem[16'h4D55] = 8'h00;
mem[16'h4D56] = 8'h72;
mem[16'h4D57] = 8'h09;
mem[16'h4D58] = 8'h72;
mem[16'h4D59] = 8'h09;
mem[16'h4D5A] = 8'h64;
mem[16'h4D5B] = 8'h04;
mem[16'h4D5C] = 8'h78;
mem[16'h4D5D] = 8'h03;
mem[16'h4D5E] = 8'h70;
mem[16'h4D5F] = 8'h01;
mem[16'h4D60] = 8'h70;
mem[16'h4D61] = 8'h01;
mem[16'h4D62] = 8'h70;
mem[16'h4D63] = 8'h01;
mem[16'h4D64] = 8'h78;
mem[16'h4D65] = 8'h03;
mem[16'h4D66] = 8'h6C;
mem[16'h4D67] = 8'h06;
mem[16'h4D68] = 8'h0C;
mem[16'h4D69] = 8'h06;
mem[16'h4D6A] = 8'h04;
mem[16'h4D6B] = 8'h04;
mem[16'h4D6C] = 8'h0A;
mem[16'h4D6D] = 8'h0A;
mem[16'h4D6E] = 8'h0A;
mem[16'h4D6F] = 8'h0A;
mem[16'h4D70] = 8'h04;
mem[16'h4D71] = 8'h04;
mem[16'h4D72] = 8'h0C;
mem[16'h4D73] = 8'h06;
mem[16'h4D74] = 8'h6C;
mem[16'h4D75] = 8'h06;
mem[16'h4D76] = 8'h78;
mem[16'h4D77] = 8'h03;
mem[16'h4D78] = 8'h70;
mem[16'h4D79] = 8'h01;
mem[16'h4D7A] = 8'h70;
mem[16'h4D7B] = 8'h01;
mem[16'h4D7C] = 8'h70;
mem[16'h4D7D] = 8'h01;
mem[16'h4D7E] = 8'h78;
mem[16'h4D7F] = 8'h03;
mem[16'h4D80] = 8'h64;
mem[16'h4D81] = 8'h04;
mem[16'h4D82] = 8'h72;
mem[16'h4D83] = 8'h09;
mem[16'h4D84] = 8'h72;
mem[16'h4D85] = 8'h09;
mem[16'h4D86] = 8'h60;
mem[16'h4D87] = 8'h00;
mem[16'h4D88] = 8'h00;
mem[16'h4D89] = 8'h00;
mem[16'h4D8A] = 8'h06;
mem[16'h4D8B] = 8'h20;
mem[16'h4D8C] = 8'h08;
mem[16'h4D8D] = 8'h1C;
mem[16'h4D8E] = 8'h10;
mem[16'h4D8F] = 8'h2E;
mem[16'h4D90] = 8'h76;
mem[16'h4D91] = 8'h03;
mem[16'h4D92] = 8'h7F;
mem[16'h4D93] = 8'h07;
mem[16'h4D94] = 8'h7F;
mem[16'h4D95] = 8'h07;
mem[16'h4D96] = 8'h76;
mem[16'h4D97] = 8'h03;
mem[16'h4D98] = 8'h10;
mem[16'h4D99] = 8'h2E;
mem[16'h4D9A] = 8'h08;
mem[16'h4D9B] = 8'h1C;
mem[16'h4D9C] = 8'h06;
mem[16'h4D9D] = 8'h20;
mem[16'h4D9E] = 8'h00;
mem[16'h4D9F] = 8'h00;
mem[16'h4DA0] = 8'h01;
mem[16'h4DA1] = 8'h18;
mem[16'h4DA2] = 8'h0E;
mem[16'h4DA3] = 8'h04;
mem[16'h4DA4] = 8'h1D;
mem[16'h4DA5] = 8'h02;
mem[16'h4DA6] = 8'h70;
mem[16'h4DA7] = 8'h1B;
mem[16'h4DA8] = 8'h78;
mem[16'h4DA9] = 8'h3F;
mem[16'h4DAA] = 8'h78;
mem[16'h4DAB] = 8'h3F;
mem[16'h4DAC] = 8'h70;
mem[16'h4DAD] = 8'h1B;
mem[16'h4DAE] = 8'h1D;
mem[16'h4DAF] = 8'h02;
mem[16'h4DB0] = 8'h0E;
mem[16'h4DB1] = 8'h04;
mem[16'h4DB2] = 8'h01;
mem[16'h4DB3] = 8'h18;
mem[16'h4DB4] = 8'hA9;
mem[16'h4DB5] = 8'h7E;
mem[16'h4DB6] = 8'h8D;
mem[16'h4DB7] = 8'hCF;
mem[16'h4DB8] = 8'h4D;
mem[16'h4DB9] = 8'hA9;
mem[16'h4DBA] = 8'hAF;
mem[16'h4DBB] = 8'h8D;
mem[16'h4DBC] = 8'hD0;
mem[16'h4DBD] = 8'h4D;
mem[16'h4DBE] = 8'hAD;
mem[16'h4DBF] = 8'h10;
mem[16'h4DC0] = 8'hC0;
mem[16'h4DC1] = 8'hA9;
mem[16'h4DC2] = 8'h00;
mem[16'h4DC3] = 8'h85;
mem[16'h4DC4] = 8'h77;
mem[16'h4DC5] = 8'h85;
mem[16'h4DC6] = 8'h87;
mem[16'h4DC7] = 8'h85;
mem[16'h4DC8] = 8'h86;
mem[16'h4DC9] = 8'h85;
mem[16'h4DCA] = 8'h88;
mem[16'h4DCB] = 8'h20;
mem[16'h4DCC] = 8'hD9;
mem[16'h4DCD] = 8'h4C;
mem[16'h4DCE] = 8'h60;
mem[16'h4DCF] = 8'h7E;
mem[16'h4DD0] = 8'hAF;
mem[16'h4DD1] = 8'hA9;
mem[16'h4DD2] = 8'h02;
mem[16'h4DD3] = 8'h8D;
mem[16'h4DD4] = 8'hAD;
mem[16'h4DD5] = 8'h4A;
mem[16'h4DD6] = 8'h8D;
mem[16'h4DD7] = 8'hB1;
mem[16'h4DD8] = 8'h4A;
mem[16'h4DD9] = 8'h8D;
mem[16'h4DDA] = 8'h63;
mem[16'h4DDB] = 8'h5E;
mem[16'h4DDC] = 8'hA9;
mem[16'h4DDD] = 8'h06;
mem[16'h4DDE] = 8'h8D;
mem[16'h4DDF] = 8'hAF;
mem[16'h4DE0] = 8'h4A;
mem[16'h4DE1] = 8'hA9;
mem[16'h4DE2] = 8'h50;
mem[16'h4DE3] = 8'h8D;
mem[16'h4DE4] = 8'hB1;
mem[16'h4DE5] = 8'h85;
mem[16'h4DE6] = 8'h8D;
mem[16'h4DE7] = 8'hB0;
mem[16'h4DE8] = 8'h85;
mem[16'h4DE9] = 8'hA9;
mem[16'h4DEA] = 8'h01;
mem[16'h4DEB] = 8'h8D;
mem[16'h4DEC] = 8'h5A;
mem[16'h4DED] = 8'h74;
mem[16'h4DEE] = 8'h8D;
mem[16'h4DEF] = 8'hB2;
mem[16'h4DF0] = 8'h4A;
mem[16'h4DF1] = 8'hA9;
mem[16'h4DF2] = 8'h03;
mem[16'h4DF3] = 8'h8D;
mem[16'h4DF4] = 8'hAA;
mem[16'h4DF5] = 8'h4A;
mem[16'h4DF6] = 8'h8D;
mem[16'h4DF7] = 8'hAE;
mem[16'h4DF8] = 8'h4A;
mem[16'h4DF9] = 8'h8D;
mem[16'h4DFA] = 8'hAB;
mem[16'h4DFB] = 8'h4A;
mem[16'h4DFC] = 8'h8D;
mem[16'h4DFD] = 8'hB3;
mem[16'h4DFE] = 8'h4A;
mem[16'h4DFF] = 8'h8D;
mem[16'h4E00] = 8'hAC;
mem[16'h4E01] = 8'h4A;
mem[16'h4E02] = 8'hA9;
mem[16'h4E03] = 8'h38;
mem[16'h4E04] = 8'h8D;
mem[16'h4E05] = 8'h4E;
mem[16'h4E06] = 8'h5E;
mem[16'h4E07] = 8'hA9;
mem[16'h4E08] = 8'h78;
mem[16'h4E09] = 8'h8D;
mem[16'h4E0A] = 8'h6B;
mem[16'h4E0B] = 8'h53;
mem[16'h4E0C] = 8'hA9;
mem[16'h4E0D] = 8'hB4;
mem[16'h4E0E] = 8'h8D;
mem[16'h4E0F] = 8'h7A;
mem[16'h4E10] = 8'h53;
mem[16'h4E11] = 8'hA9;
mem[16'h4E12] = 8'hF0;
mem[16'h4E13] = 8'h8D;
mem[16'h4E14] = 8'hD1;
mem[16'h4E15] = 8'h4F;
mem[16'h4E16] = 8'hA9;
mem[16'h4E17] = 8'h40;
mem[16'h4E18] = 8'h8D;
mem[16'h4E19] = 8'hBD;
mem[16'h4E1A] = 8'h5F;
mem[16'h4E1B] = 8'hA9;
mem[16'h4E1C] = 8'h50;
mem[16'h4E1D] = 8'h8D;
mem[16'h4E1E] = 8'hF8;
mem[16'h4E1F] = 8'h5D;
mem[16'h4E20] = 8'hA9;
mem[16'h4E21] = 8'h78;
mem[16'h4E22] = 8'h8D;
mem[16'h4E23] = 8'h5E;
mem[16'h4E24] = 8'h5F;
mem[16'h4E25] = 8'hA9;
mem[16'h4E26] = 8'h54;
mem[16'h4E27] = 8'h8D;
mem[16'h4E28] = 8'hCA;
mem[16'h4E29] = 8'h5D;
mem[16'h4E2A] = 8'hA9;
mem[16'h4E2B] = 8'hA0;
mem[16'h4E2C] = 8'h8D;
mem[16'h4E2D] = 8'h1F;
mem[16'h4E2E] = 8'h51;
mem[16'h4E2F] = 8'hA9;
mem[16'h4E30] = 8'h30;
mem[16'h4E31] = 8'h8D;
mem[16'h4E32] = 8'h27;
mem[16'h4E33] = 8'h53;
mem[16'h4E34] = 8'hA9;
mem[16'h4E35] = 8'h1E;
mem[16'h4E36] = 8'h8D;
mem[16'h4E37] = 8'hDD;
mem[16'h4E38] = 8'h91;
mem[16'h4E39] = 8'h8D;
mem[16'h4E3A] = 8'hDC;
mem[16'h4E3B] = 8'h91;
mem[16'h4E3C] = 8'hA9;
mem[16'h4E3D] = 8'hC8;
mem[16'h4E3E] = 8'h8D;
mem[16'h4E3F] = 8'h22;
mem[16'h4E40] = 8'h43;
mem[16'h4E41] = 8'hA9;
mem[16'h4E42] = 8'hB4;
mem[16'h4E43] = 8'h8D;
mem[16'h4E44] = 8'h57;
mem[16'h4E45] = 8'h42;
mem[16'h4E46] = 8'h20;
mem[16'h4E47] = 8'h79;
mem[16'h4E48] = 8'h4A;
mem[16'h4E49] = 8'hA9;
mem[16'h4E4A] = 8'h54;
mem[16'h4E4B] = 8'h85;
mem[16'h4E4C] = 8'h5E;
mem[16'h4E4D] = 8'hA9;
mem[16'h4E4E] = 8'h4E;
mem[16'h4E4F] = 8'h85;
mem[16'h4E50] = 8'h5F;
mem[16'h4E51] = 8'h4C;
mem[16'h4E52] = 8'h18;
mem[16'h4E53] = 8'h40;
mem[16'h4E54] = 8'hA9;
mem[16'h4E55] = 8'h64;
mem[16'h4E56] = 8'h8D;
mem[16'h4E57] = 8'hB0;
mem[16'h4E58] = 8'h85;
mem[16'h4E59] = 8'h8D;
mem[16'h4E5A] = 8'hB1;
mem[16'h4E5B] = 8'h85;
mem[16'h4E5C] = 8'hA9;
mem[16'h4E5D] = 8'h02;
mem[16'h4E5E] = 8'h8D;
mem[16'h4E5F] = 8'hB1;
mem[16'h4E60] = 8'h4A;
mem[16'h4E61] = 8'hA9;
mem[16'h4E62] = 8'h01;
mem[16'h4E63] = 8'h8D;
mem[16'h4E64] = 8'h5A;
mem[16'h4E65] = 8'h74;
mem[16'h4E66] = 8'hA9;
mem[16'h4E67] = 8'h03;
mem[16'h4E68] = 8'h8D;
mem[16'h4E69] = 8'hB3;
mem[16'h4E6A] = 8'h4A;
mem[16'h4E6B] = 8'h8D;
mem[16'h4E6C] = 8'hAE;
mem[16'h4E6D] = 8'h4A;
mem[16'h4E6E] = 8'h8D;
mem[16'h4E6F] = 8'hAD;
mem[16'h4E70] = 8'h4A;
mem[16'h4E71] = 8'h8D;
mem[16'h4E72] = 8'hAB;
mem[16'h4E73] = 8'h4A;
mem[16'h4E74] = 8'h8D;
mem[16'h4E75] = 8'hAA;
mem[16'h4E76] = 8'h4A;
mem[16'h4E77] = 8'hA9;
mem[16'h4E78] = 8'h04;
mem[16'h4E79] = 8'h8D;
mem[16'h4E7A] = 8'hAC;
mem[16'h4E7B] = 8'h4A;
mem[16'h4E7C] = 8'h8D;
mem[16'h4E7D] = 8'hAF;
mem[16'h4E7E] = 8'h4A;
mem[16'h4E7F] = 8'hA9;
mem[16'h4E80] = 8'h66;
mem[16'h4E81] = 8'h8D;
mem[16'h4E82] = 8'h4E;
mem[16'h4E83] = 8'h5E;
mem[16'h4E84] = 8'hA9;
mem[16'h4E85] = 8'h64;
mem[16'h4E86] = 8'h8D;
mem[16'h4E87] = 8'hE3;
mem[16'h4E88] = 8'h51;
mem[16'h4E89] = 8'hA9;
mem[16'h4E8A] = 8'hC8;
mem[16'h4E8B] = 8'h8D;
mem[16'h4E8C] = 8'hF2;
mem[16'h4E8D] = 8'h51;
mem[16'h4E8E] = 8'hA9;
mem[16'h4E8F] = 8'h1C;
mem[16'h4E90] = 8'h8D;
mem[16'h4E91] = 8'hDD;
mem[16'h4E92] = 8'h91;
mem[16'h4E93] = 8'hA9;
mem[16'h4E94] = 8'h54;
mem[16'h4E95] = 8'h8D;
mem[16'h4E96] = 8'h5E;
mem[16'h4E97] = 8'h5F;
mem[16'h4E98] = 8'hA9;
mem[16'h4E99] = 8'h24;
mem[16'h4E9A] = 8'h8D;
mem[16'h4E9B] = 8'h27;
mem[16'h4E9C] = 8'h53;
mem[16'h4E9D] = 8'hA9;
mem[16'h4E9E] = 8'h10;
mem[16'h4E9F] = 8'h8D;
mem[16'h4EA0] = 8'hDF;
mem[16'h4EA1] = 8'h91;
mem[16'h4EA2] = 8'hA9;
mem[16'h4EA3] = 8'h15;
mem[16'h4EA4] = 8'h8D;
mem[16'h4EA5] = 8'hDE;
mem[16'h4EA6] = 8'h91;
mem[16'h4EA7] = 8'hA0;
mem[16'h4EA8] = 8'h01;
mem[16'h4EA9] = 8'hAD;
mem[16'h4EAA] = 8'hCE;
mem[16'h4EAB] = 8'h44;
mem[16'h4EAC] = 8'hC9;
mem[16'h4EAD] = 8'h06;
mem[16'h4EAE] = 8'h90;
mem[16'h4EAF] = 8'h02;
mem[16'h4EB0] = 8'hA0;
mem[16'h4EB1] = 8'h02;
mem[16'h4EB2] = 8'h8C;
mem[16'h4EB3] = 8'hC7;
mem[16'h4EB4] = 8'h77;
mem[16'h4EB5] = 8'hA9;
mem[16'h4EB6] = 8'h40;
mem[16'h4EB7] = 8'h8D;
mem[16'h4EB8] = 8'h0C;
mem[16'h4EB9] = 8'h54;
mem[16'h4EBA] = 8'hA9;
mem[16'h4EBB] = 8'hC8;
mem[16'h4EBC] = 8'h8D;
mem[16'h4EBD] = 8'h22;
mem[16'h4EBE] = 8'h43;
mem[16'h4EBF] = 8'hA9;
mem[16'h4EC0] = 8'hB4;
mem[16'h4EC1] = 8'h8D;
mem[16'h4EC2] = 8'h57;
mem[16'h4EC3] = 8'h42;
mem[16'h4EC4] = 8'h20;
mem[16'h4EC5] = 8'h79;
mem[16'h4EC6] = 8'h4A;
mem[16'h4EC7] = 8'hA9;
mem[16'h4EC8] = 8'hD2;
mem[16'h4EC9] = 8'h85;
mem[16'h4ECA] = 8'h5E;
mem[16'h4ECB] = 8'hA9;
mem[16'h4ECC] = 8'h4E;
mem[16'h4ECD] = 8'h85;
mem[16'h4ECE] = 8'h5F;
mem[16'h4ECF] = 8'h4C;
mem[16'h4ED0] = 8'h18;
mem[16'h4ED1] = 8'h40;
mem[16'h4ED2] = 8'hA9;
mem[16'h4ED3] = 8'h64;
mem[16'h4ED4] = 8'h8D;
mem[16'h4ED5] = 8'hB0;
mem[16'h4ED6] = 8'h85;
mem[16'h4ED7] = 8'h8D;
mem[16'h4ED8] = 8'hB1;
mem[16'h4ED9] = 8'h85;
mem[16'h4EDA] = 8'hA9;
mem[16'h4EDB] = 8'h01;
mem[16'h4EDC] = 8'h8D;
mem[16'h4EDD] = 8'h5A;
mem[16'h4EDE] = 8'h74;
mem[16'h4EDF] = 8'hA9;
mem[16'h4EE0] = 8'h02;
mem[16'h4EE1] = 8'h8D;
mem[16'h4EE2] = 8'hB1;
mem[16'h4EE3] = 8'h4A;
mem[16'h4EE4] = 8'h8D;
mem[16'h4EE5] = 8'hB3;
mem[16'h4EE6] = 8'h4A;
mem[16'h4EE7] = 8'hA9;
mem[16'h4EE8] = 8'h04;
mem[16'h4EE9] = 8'h8D;
mem[16'h4EEA] = 8'hAD;
mem[16'h4EEB] = 8'h4A;
mem[16'h4EEC] = 8'hA9;
mem[16'h4EED] = 8'h0A;
mem[16'h4EEE] = 8'h8D;
mem[16'h4EEF] = 8'hDF;
mem[16'h4EF0] = 8'h91;
mem[16'h4EF1] = 8'hA9;
mem[16'h4EF2] = 8'h14;
mem[16'h4EF3] = 8'h8D;
mem[16'h4EF4] = 8'hDD;
mem[16'h4EF5] = 8'h91;
mem[16'h4EF6] = 8'hA9;
mem[16'h4EF7] = 8'h0B;
mem[16'h4EF8] = 8'h8D;
mem[16'h4EF9] = 8'hDE;
mem[16'h4EFA] = 8'h91;
mem[16'h4EFB] = 8'hA9;
mem[16'h4EFC] = 8'h32;
mem[16'h4EFD] = 8'h8D;
mem[16'h4EFE] = 8'h27;
mem[16'h4EFF] = 8'h53;
mem[16'h4F00] = 8'hA9;
mem[16'h4F01] = 8'h40;
mem[16'h4F02] = 8'h8D;
mem[16'h4F03] = 8'h5E;
mem[16'h4F04] = 8'h5F;
mem[16'h4F05] = 8'hA9;
mem[16'h4F06] = 8'h44;
mem[16'h4F07] = 8'h8D;
mem[16'h4F08] = 8'hAF;
mem[16'h4F09] = 8'h5E;
mem[16'h4F0A] = 8'hA9;
mem[16'h4F0B] = 8'h54;
mem[16'h4F0C] = 8'h8D;
mem[16'h4F0D] = 8'hCA;
mem[16'h4F0E] = 8'h5D;
mem[16'h4F0F] = 8'hA9;
mem[16'h4F10] = 8'h8C;
mem[16'h4F11] = 8'h8D;
mem[16'h4F12] = 8'hE3;
mem[16'h4F13] = 8'h51;
mem[16'h4F14] = 8'hA9;
mem[16'h4F15] = 8'hB4;
mem[16'h4F16] = 8'h8D;
mem[16'h4F17] = 8'h57;
mem[16'h4F18] = 8'h42;
mem[16'h4F19] = 8'hA9;
mem[16'h4F1A] = 8'hC8;
mem[16'h4F1B] = 8'h8D;
mem[16'h4F1C] = 8'h22;
mem[16'h4F1D] = 8'h43;
mem[16'h4F1E] = 8'h20;
mem[16'h4F1F] = 8'h79;
mem[16'h4F20] = 8'h4A;
mem[16'h4F21] = 8'hA9;
mem[16'h4F22] = 8'h2C;
mem[16'h4F23] = 8'h85;
mem[16'h4F24] = 8'h5E;
mem[16'h4F25] = 8'hA9;
mem[16'h4F26] = 8'h4F;
mem[16'h4F27] = 8'h85;
mem[16'h4F28] = 8'h5F;
mem[16'h4F29] = 8'h4C;
mem[16'h4F2A] = 8'h18;
mem[16'h4F2B] = 8'h40;
mem[16'h4F2C] = 8'hA9;
mem[16'h4F2D] = 8'h00;
mem[16'h4F2E] = 8'h8D;
mem[16'h4F2F] = 8'hB1;
mem[16'h4F30] = 8'h4A;
mem[16'h4F31] = 8'hA9;
mem[16'h4F32] = 8'h64;
mem[16'h4F33] = 8'h8D;
mem[16'h4F34] = 8'hB0;
mem[16'h4F35] = 8'h85;
mem[16'h4F36] = 8'h8D;
mem[16'h4F37] = 8'hB1;
mem[16'h4F38] = 8'h85;
mem[16'h4F39] = 8'hA9;
mem[16'h4F3A] = 8'h01;
mem[16'h4F3B] = 8'h8D;
mem[16'h4F3C] = 8'h5A;
mem[16'h4F3D] = 8'h74;
mem[16'h4F3E] = 8'hA9;
mem[16'h4F3F] = 8'h02;
mem[16'h4F40] = 8'h8D;
mem[16'h4F41] = 8'hB3;
mem[16'h4F42] = 8'h4A;
mem[16'h4F43] = 8'hA9;
mem[16'h4F44] = 8'h04;
mem[16'h4F45] = 8'h8D;
mem[16'h4F46] = 8'hAA;
mem[16'h4F47] = 8'h4A;
mem[16'h4F48] = 8'hA9;
mem[16'h4F49] = 8'h0B;
mem[16'h4F4A] = 8'h8D;
mem[16'h4F4B] = 8'hB0;
mem[16'h4F4C] = 8'h4A;
mem[16'h4F4D] = 8'hA9;
mem[16'h4F4E] = 8'h04;
mem[16'h4F4F] = 8'h8D;
mem[16'h4F50] = 8'hAF;
mem[16'h4F51] = 8'h4A;
mem[16'h4F52] = 8'hA9;
mem[16'h4F53] = 8'h40;
mem[16'h4F54] = 8'h8D;
mem[16'h4F55] = 8'h8F;
mem[16'h4F56] = 8'h5F;
mem[16'h4F57] = 8'hA9;
mem[16'h4F58] = 8'hB4;
mem[16'h4F59] = 8'h8D;
mem[16'h4F5A] = 8'hE3;
mem[16'h4F5B] = 8'h51;
mem[16'h4F5C] = 8'hA9;
mem[16'h4F5D] = 8'h52;
mem[16'h4F5E] = 8'h8D;
mem[16'h4F5F] = 8'hAF;
mem[16'h4F60] = 8'h5E;
mem[16'h4F61] = 8'h20;
mem[16'h4F62] = 8'h79;
mem[16'h4F63] = 8'h4A;
mem[16'h4F64] = 8'hA9;
mem[16'h4F65] = 8'h55;
mem[16'h4F66] = 8'h85;
mem[16'h4F67] = 8'h5E;
mem[16'h4F68] = 8'hA9;
mem[16'h4F69] = 8'h49;
mem[16'h4F6A] = 8'h85;
mem[16'h4F6B] = 8'h5F;
mem[16'h4F6C] = 8'h4C;
mem[16'h4F6D] = 8'h18;
mem[16'h4F6E] = 8'h40;
mem[16'h4F6F] = 8'h20;
mem[16'h4F70] = 8'h05;
mem[16'h4F71] = 8'h08;
mem[16'h4F72] = 8'h10;
mem[16'h4F73] = 8'h00;
mem[16'h4F74] = 8'h00;
mem[16'h4F75] = 8'h62;
mem[16'h4F76] = 8'h47;
mem[16'h4F77] = 8'h72;
mem[16'h4F78] = 8'h4F;
mem[16'h4F79] = 8'h72;
mem[16'h4F7A] = 8'h4F;
mem[16'h4F7B] = 8'h72;
mem[16'h4F7C] = 8'h4F;
mem[16'h4F7D] = 8'h62;
mem[16'h4F7E] = 8'h47;
mem[16'h4F7F] = 8'h00;
mem[16'h4F80] = 8'h00;
mem[16'h4F81] = 8'h08;
mem[16'h4F82] = 8'h10;
mem[16'h4F83] = 8'h20;
mem[16'h4F84] = 8'h05;
mem[16'h4F85] = 8'h00;
mem[16'h4F86] = 8'h00;
mem[16'h4F87] = 8'h00;
mem[16'h4F88] = 8'h00;
mem[16'h4F89] = 8'h20;
mem[16'h4F8A] = 8'h05;
mem[16'h4F8B] = 8'h00;
mem[16'h4F8C] = 8'h00;
mem[16'h4F8D] = 8'h48;
mem[16'h4F8E] = 8'h13;
mem[16'h4F8F] = 8'h68;
mem[16'h4F90] = 8'h17;
mem[16'h4F91] = 8'h48;
mem[16'h4F92] = 8'h13;
mem[16'h4F93] = 8'h00;
mem[16'h4F94] = 8'h00;
mem[16'h4F95] = 8'h20;
mem[16'h4F96] = 8'h05;
mem[16'h4F97] = 8'hA9;
mem[16'h4F98] = 8'h00;
mem[16'h4F99] = 8'h8D;
mem[16'h4F9A] = 8'hF8;
mem[16'h4F9B] = 8'h4F;
mem[16'h4F9C] = 8'h8D;
mem[16'h4F9D] = 8'h19;
mem[16'h4F9E] = 8'h51;
mem[16'h4F9F] = 8'h8D;
mem[16'h4FA0] = 8'h1A;
mem[16'h4FA1] = 8'h51;
mem[16'h4FA2] = 8'h8D;
mem[16'h4FA3] = 8'h1B;
mem[16'h4FA4] = 8'h51;
mem[16'h4FA5] = 8'h8D;
mem[16'h4FA6] = 8'h1C;
mem[16'h4FA7] = 8'h51;
mem[16'h4FA8] = 8'h8D;
mem[16'h4FA9] = 8'h1D;
mem[16'h4FAA] = 8'h51;
mem[16'h4FAB] = 8'h8D;
mem[16'h4FAC] = 8'h1E;
mem[16'h4FAD] = 8'h51;
mem[16'h4FAE] = 8'hA9;
mem[16'h4FAF] = 8'h01;
mem[16'h4FB0] = 8'h8D;
mem[16'h4FB1] = 8'h10;
mem[16'h4FB2] = 8'h51;
mem[16'h4FB3] = 8'h8D;
mem[16'h4FB4] = 8'h11;
mem[16'h4FB5] = 8'h51;
mem[16'h4FB6] = 8'h8D;
mem[16'h4FB7] = 8'h12;
mem[16'h4FB8] = 8'h51;
mem[16'h4FB9] = 8'hAD;
mem[16'h4FBA] = 8'h1F;
mem[16'h4FBB] = 8'h51;
mem[16'h4FBC] = 8'h8D;
mem[16'h4FBD] = 8'h16;
mem[16'h4FBE] = 8'h51;
mem[16'h4FBF] = 8'h8D;
mem[16'h4FC0] = 8'h17;
mem[16'h4FC1] = 8'h51;
mem[16'h4FC2] = 8'h8D;
mem[16'h4FC3] = 8'h18;
mem[16'h4FC4] = 8'h51;
mem[16'h4FC5] = 8'hA9;
mem[16'h4FC6] = 8'h01;
mem[16'h4FC7] = 8'h8D;
mem[16'h4FC8] = 8'hF8;
mem[16'h4FC9] = 8'h4F;
mem[16'h4FCA] = 8'h20;
mem[16'h4FCB] = 8'hF7;
mem[16'h4FCC] = 8'h4F;
mem[16'h4FCD] = 8'hAD;
mem[16'h4FCE] = 8'h10;
mem[16'h4FCF] = 8'h51;
mem[16'h4FD0] = 8'hC9;
mem[16'h4FD1] = 8'hAA;
mem[16'h4FD2] = 8'h90;
mem[16'h4FD3] = 8'hF6;
mem[16'h4FD4] = 8'hA9;
mem[16'h4FD5] = 8'h02;
mem[16'h4FD6] = 8'hCD;
mem[16'h4FD7] = 8'hB2;
mem[16'h4FD8] = 8'h4A;
mem[16'h4FD9] = 8'hF0;
mem[16'h4FDA] = 8'h02;
mem[16'h4FDB] = 8'hB0;
mem[16'h4FDC] = 8'h19;
mem[16'h4FDD] = 8'h8D;
mem[16'h4FDE] = 8'hF8;
mem[16'h4FDF] = 8'h4F;
mem[16'h4FE0] = 8'h20;
mem[16'h4FE1] = 8'hF7;
mem[16'h4FE2] = 8'h4F;
mem[16'h4FE3] = 8'hAD;
mem[16'h4FE4] = 8'h10;
mem[16'h4FE5] = 8'h51;
mem[16'h4FE6] = 8'hC9;
mem[16'h4FE7] = 8'hB0;
mem[16'h4FE8] = 8'h90;
mem[16'h4FE9] = 8'hF6;
mem[16'h4FEA] = 8'hA9;
mem[16'h4FEB] = 8'h03;
mem[16'h4FEC] = 8'hCD;
mem[16'h4FED] = 8'hB2;
mem[16'h4FEE] = 8'h4A;
mem[16'h4FEF] = 8'hF0;
mem[16'h4FF0] = 8'h02;
mem[16'h4FF1] = 8'hB0;
mem[16'h4FF2] = 8'h03;
mem[16'h4FF3] = 8'h8D;
mem[16'h4FF4] = 8'hF8;
mem[16'h4FF5] = 8'h4F;
mem[16'h4FF6] = 8'h60;
mem[16'h4FF7] = 8'hA2;
mem[16'h4FF8] = 8'h02;
mem[16'h4FF9] = 8'hCA;
mem[16'h4FFA] = 8'h30;
mem[16'h4FFB] = 8'h62;
mem[16'h4FFC] = 8'h86;
mem[16'h4FFD] = 8'h70;
mem[16'h4FFE] = 8'h20;
mem[16'h4FFF] = 8'hD2;
mem[16'h5000] = 8'h50;
mem[16'h5001] = 8'hA6;
mem[16'h5002] = 8'h70;
mem[16'h5003] = 8'hBD;
mem[16'h5004] = 8'h10;
mem[16'h5005] = 8'h51;
mem[16'h5006] = 8'hAC;
mem[16'h5007] = 8'hB2;
mem[16'h5008] = 8'h4A;
mem[16'h5009] = 8'hC0;
mem[16'h500A] = 8'h01;
mem[16'h500B] = 8'hF0;
mem[16'h500C] = 8'h04;
mem[16'h500D] = 8'hC9;
mem[16'h500E] = 8'hFC;
mem[16'h500F] = 8'hB0;
mem[16'h5010] = 8'h2A;
mem[16'h5011] = 8'h18;
mem[16'h5012] = 8'h69;
mem[16'h5013] = 8'h04;
mem[16'h5014] = 8'h9D;
mem[16'h5015] = 8'h10;
mem[16'h5016] = 8'h51;
mem[16'h5017] = 8'h20;
mem[16'h5018] = 8'h81;
mem[16'h5019] = 8'h50;
mem[16'h501A] = 8'hA6;
mem[16'h501B] = 8'h70;
mem[16'h501C] = 8'hAC;
mem[16'h501D] = 8'hB2;
mem[16'h501E] = 8'h4A;
mem[16'h501F] = 8'hC0;
mem[16'h5020] = 8'h01;
mem[16'h5021] = 8'hD0;
mem[16'h5022] = 8'hD6;
mem[16'h5023] = 8'hBD;
mem[16'h5024] = 8'h10;
mem[16'h5025] = 8'h51;
mem[16'h5026] = 8'h38;
mem[16'h5027] = 8'hFD;
mem[16'h5028] = 8'h16;
mem[16'h5029] = 8'h51;
mem[16'h502A] = 8'hC9;
mem[16'h502B] = 8'hFD;
mem[16'h502C] = 8'h90;
mem[16'h502D] = 8'hCB;
mem[16'h502E] = 8'h20;
mem[16'h502F] = 8'hB1;
mem[16'h5030] = 8'h50;
mem[16'h5031] = 8'hA6;
mem[16'h5032] = 8'h70;
mem[16'h5033] = 8'hA9;
mem[16'h5034] = 8'h00;
mem[16'h5035] = 8'h9D;
mem[16'h5036] = 8'h19;
mem[16'h5037] = 8'h51;
mem[16'h5038] = 8'h4C;
mem[16'h5039] = 8'hF9;
mem[16'h503A] = 8'h4F;
mem[16'h503B] = 8'hBD;
mem[16'h503C] = 8'h16;
mem[16'h503D] = 8'h51;
mem[16'h503E] = 8'h38;
mem[16'h503F] = 8'hE9;
mem[16'h5040] = 8'h04;
mem[16'h5041] = 8'h9D;
mem[16'h5042] = 8'h16;
mem[16'h5043] = 8'h51;
mem[16'h5044] = 8'hD0;
mem[16'h5045] = 8'hB3;
mem[16'h5046] = 8'h20;
mem[16'h5047] = 8'h88;
mem[16'h5048] = 8'h50;
mem[16'h5049] = 8'hA6;
mem[16'h504A] = 8'h70;
mem[16'h504B] = 8'hA9;
mem[16'h504C] = 8'h00;
mem[16'h504D] = 8'h9D;
mem[16'h504E] = 8'h19;
mem[16'h504F] = 8'h51;
mem[16'h5050] = 8'hA9;
mem[16'h5051] = 8'h01;
mem[16'h5052] = 8'h9D;
mem[16'h5053] = 8'h10;
mem[16'h5054] = 8'h51;
mem[16'h5055] = 8'hAD;
mem[16'h5056] = 8'h1F;
mem[16'h5057] = 8'h51;
mem[16'h5058] = 8'h9D;
mem[16'h5059] = 8'h16;
mem[16'h505A] = 8'h51;
mem[16'h505B] = 8'h4C;
mem[16'h505C] = 8'hF9;
mem[16'h505D] = 8'h4F;
mem[16'h505E] = 8'h60;
mem[16'h505F] = 8'hA9;
mem[16'h5060] = 8'h12;
mem[16'h5061] = 8'h8D;
mem[16'h5062] = 8'h24;
mem[16'h5063] = 8'h8C;
mem[16'h5064] = 8'hA9;
mem[16'h5065] = 8'h6F;
mem[16'h5066] = 8'hA0;
mem[16'h5067] = 8'h50;
mem[16'h5068] = 8'h20;
mem[16'h5069] = 8'h2B;
mem[16'h506A] = 8'h8C;
mem[16'h506B] = 8'h20;
mem[16'h506C] = 8'hA8;
mem[16'h506D] = 8'h8B;
mem[16'h506E] = 8'h60;
mem[16'h506F] = 8'h70;
mem[16'h5070] = 8'h01;
mem[16'h5071] = 8'h3C;
mem[16'h5072] = 8'h00;
mem[16'h5073] = 8'h0F;
mem[16'h5074] = 8'h00;
mem[16'h5075] = 8'h0F;
mem[16'h5076] = 8'h00;
mem[16'h5077] = 8'h0F;
mem[16'h5078] = 8'h00;
mem[16'h5079] = 8'h0F;
mem[16'h507A] = 8'h00;
mem[16'h507B] = 8'h0F;
mem[16'h507C] = 8'h00;
mem[16'h507D] = 8'h3C;
mem[16'h507E] = 8'h00;
mem[16'h507F] = 8'h70;
mem[16'h5080] = 8'h01;
mem[16'h5081] = 8'hA6;
mem[16'h5082] = 8'h70;
mem[16'h5083] = 8'hBD;
mem[16'h5084] = 8'h19;
mem[16'h5085] = 8'h51;
mem[16'h5086] = 8'hD0;
mem[16'h5087] = 8'h28;
mem[16'h5088] = 8'hA6;
mem[16'h5089] = 8'h70;
mem[16'h508A] = 8'hBD;
mem[16'h508B] = 8'h13;
mem[16'h508C] = 8'h51;
mem[16'h508D] = 8'h85;
mem[16'h508E] = 8'h56;
mem[16'h508F] = 8'hBD;
mem[16'h5090] = 8'h10;
mem[16'h5091] = 8'h51;
mem[16'h5092] = 8'h38;
mem[16'h5093] = 8'hFD;
mem[16'h5094] = 8'h16;
mem[16'h5095] = 8'h51;
mem[16'h5096] = 8'h90;
mem[16'h5097] = 8'h18;
mem[16'h5098] = 8'h85;
mem[16'h5099] = 8'h57;
mem[16'h509A] = 8'hA9;
mem[16'h509B] = 8'h09;
mem[16'h509C] = 8'h8D;
mem[16'h509D] = 8'hC0;
mem[16'h509E] = 8'h65;
mem[16'h509F] = 8'hA9;
mem[16'h50A0] = 8'hC9;
mem[16'h50A1] = 8'hA0;
mem[16'h50A2] = 8'h50;
mem[16'h50A3] = 8'h20;
mem[16'h50A4] = 8'hC7;
mem[16'h50A5] = 8'h65;
mem[16'h50A6] = 8'h20;
mem[16'h50A7] = 8'h6A;
mem[16'h50A8] = 8'h65;
mem[16'h50A9] = 8'hA6;
mem[16'h50AA] = 8'h70;
mem[16'h50AB] = 8'hA9;
mem[16'h50AC] = 8'h01;
mem[16'h50AD] = 8'h9D;
mem[16'h50AE] = 8'h19;
mem[16'h50AF] = 8'h51;
mem[16'h50B0] = 8'h60;
mem[16'h50B1] = 8'hA6;
mem[16'h50B2] = 8'h70;
mem[16'h50B3] = 8'hBD;
mem[16'h50B4] = 8'h19;
mem[16'h50B5] = 8'h51;
mem[16'h50B6] = 8'hF0;
mem[16'h50B7] = 8'hF8;
mem[16'h50B8] = 8'hBD;
mem[16'h50B9] = 8'h13;
mem[16'h50BA] = 8'h51;
mem[16'h50BB] = 8'h85;
mem[16'h50BC] = 8'h56;
mem[16'h50BD] = 8'hBD;
mem[16'h50BE] = 8'h10;
mem[16'h50BF] = 8'h51;
mem[16'h50C0] = 8'h38;
mem[16'h50C1] = 8'hFD;
mem[16'h50C2] = 8'h16;
mem[16'h50C3] = 8'h51;
mem[16'h50C4] = 8'h85;
mem[16'h50C5] = 8'h57;
mem[16'h50C6] = 8'h4C;
mem[16'h50C7] = 8'h9A;
mem[16'h50C8] = 8'h50;
mem[16'h50C9] = 8'h0F;
mem[16'h50CA] = 8'h03;
mem[16'h50CB] = 8'h00;
mem[16'h50CC] = 8'h00;
mem[16'h50CD] = 8'h00;
mem[16'h50CE] = 8'h00;
mem[16'h50CF] = 8'h00;
mem[16'h50D0] = 8'h03;
mem[16'h50D1] = 8'h0F;
mem[16'h50D2] = 8'hA6;
mem[16'h50D3] = 8'h70;
mem[16'h50D4] = 8'hBD;
mem[16'h50D5] = 8'h13;
mem[16'h50D6] = 8'h51;
mem[16'h50D7] = 8'h85;
mem[16'h50D8] = 8'h56;
mem[16'h50D9] = 8'h85;
mem[16'h50DA] = 8'h6F;
mem[16'h50DB] = 8'hBD;
mem[16'h50DC] = 8'h10;
mem[16'h50DD] = 8'h51;
mem[16'h50DE] = 8'h85;
mem[16'h50DF] = 8'h57;
mem[16'h50E0] = 8'hC9;
mem[16'h50E1] = 8'hFD;
mem[16'h50E2] = 8'hF0;
mem[16'h50E3] = 8'h08;
mem[16'h50E4] = 8'hB0;
mem[16'h50E5] = 8'h09;
mem[16'h50E6] = 8'h20;
mem[16'h50E7] = 8'h20;
mem[16'h50E8] = 8'h51;
mem[16'h50E9] = 8'h4C;
mem[16'h50EA] = 8'hEF;
mem[16'h50EB] = 8'h50;
mem[16'h50EC] = 8'h20;
mem[16'h50ED] = 8'h5D;
mem[16'h50EE] = 8'h51;
mem[16'h50EF] = 8'hA6;
mem[16'h50F0] = 8'h70;
mem[16'h50F1] = 8'hA5;
mem[16'h50F2] = 8'h57;
mem[16'h50F3] = 8'h38;
mem[16'h50F4] = 8'hFD;
mem[16'h50F5] = 8'h16;
mem[16'h50F6] = 8'h51;
mem[16'h50F7] = 8'h90;
mem[16'h50F8] = 8'h0A;
mem[16'h50F9] = 8'h85;
mem[16'h50FA] = 8'h57;
mem[16'h50FB] = 8'hA5;
mem[16'h50FC] = 8'h6F;
mem[16'h50FD] = 8'h85;
mem[16'h50FE] = 8'h56;
mem[16'h50FF] = 8'h20;
mem[16'h5100] = 8'h5F;
mem[16'h5101] = 8'h50;
mem[16'h5102] = 8'h60;
mem[16'h5103] = 8'hAC;
mem[16'h5104] = 8'hB2;
mem[16'h5105] = 8'h4A;
mem[16'h5106] = 8'hC0;
mem[16'h5107] = 8'h01;
mem[16'h5108] = 8'hD0;
mem[16'h5109] = 8'h05;
mem[16'h510A] = 8'hBC;
mem[16'h510B] = 8'h19;
mem[16'h510C] = 8'h51;
mem[16'h510D] = 8'hD0;
mem[16'h510E] = 8'hEA;
mem[16'h510F] = 8'h60;
mem[16'h5110] = 8'hB1;
mem[16'h5111] = 8'h05;
mem[16'h5112] = 8'h01;
mem[16'h5113] = 8'h33;
mem[16'h5114] = 8'h33;
mem[16'h5115] = 8'h33;
mem[16'h5116] = 8'h64;
mem[16'h5117] = 8'h64;
mem[16'h5118] = 8'h64;
mem[16'h5119] = 8'h01;
mem[16'h511A] = 8'h00;
mem[16'h511B] = 8'h00;
mem[16'h511C] = 8'h09;
mem[16'h511D] = 8'h09;
mem[16'h511E] = 8'h00;
mem[16'h511F] = 8'h64;
mem[16'h5120] = 8'hBD;
mem[16'h5121] = 8'h1C;
mem[16'h5122] = 8'h51;
mem[16'h5123] = 8'hD0;
mem[16'h5124] = 8'h12;
mem[16'h5125] = 8'hA9;
mem[16'h5126] = 8'h79;
mem[16'h5127] = 8'hA0;
mem[16'h5128] = 8'h51;
mem[16'h5129] = 8'h20;
mem[16'h512A] = 8'hC7;
mem[16'h512B] = 8'h65;
mem[16'h512C] = 8'hA9;
mem[16'h512D] = 8'h09;
mem[16'h512E] = 8'h8D;
mem[16'h512F] = 8'hC0;
mem[16'h5130] = 8'h65;
mem[16'h5131] = 8'h9D;
mem[16'h5132] = 8'h1C;
mem[16'h5133] = 8'h51;
mem[16'h5134] = 8'h20;
mem[16'h5135] = 8'h6A;
mem[16'h5136] = 8'h65;
mem[16'h5137] = 8'hA6;
mem[16'h5138] = 8'h70;
mem[16'h5139] = 8'hBD;
mem[16'h513A] = 8'h13;
mem[16'h513B] = 8'h51;
mem[16'h513C] = 8'h85;
mem[16'h513D] = 8'h56;
mem[16'h513E] = 8'hBC;
mem[16'h513F] = 8'h10;
mem[16'h5140] = 8'h51;
mem[16'h5141] = 8'h84;
mem[16'h5142] = 8'h57;
mem[16'h5143] = 8'hB9;
mem[16'h5144] = 8'h3E;
mem[16'h5145] = 8'h8C;
mem[16'h5146] = 8'hAA;
mem[16'h5147] = 8'hBD;
mem[16'h5148] = 8'h94;
mem[16'h5149] = 8'h8E;
mem[16'h514A] = 8'hAA;
mem[16'h514B] = 8'hBD;
mem[16'h514C] = 8'h74;
mem[16'h514D] = 8'h62;
mem[16'h514E] = 8'hBC;
mem[16'h514F] = 8'h7B;
mem[16'h5150] = 8'h62;
mem[16'h5151] = 8'h20;
mem[16'h5152] = 8'h3B;
mem[16'h5153] = 8'h8B;
mem[16'h5154] = 8'hA9;
mem[16'h5155] = 8'h1B;
mem[16'h5156] = 8'h8D;
mem[16'h5157] = 8'h34;
mem[16'h5158] = 8'h8B;
mem[16'h5159] = 8'h20;
mem[16'h515A] = 8'hF0;
mem[16'h515B] = 8'h8A;
mem[16'h515C] = 8'h60;
mem[16'h515D] = 8'hBD;
mem[16'h515E] = 8'h1C;
mem[16'h515F] = 8'h51;
mem[16'h5160] = 8'hF0;
mem[16'h5161] = 8'h16;
mem[16'h5162] = 8'hA9;
mem[16'h5163] = 8'h79;
mem[16'h5164] = 8'hA0;
mem[16'h5165] = 8'h51;
mem[16'h5166] = 8'h20;
mem[16'h5167] = 8'hC7;
mem[16'h5168] = 8'h65;
mem[16'h5169] = 8'hA9;
mem[16'h516A] = 8'h09;
mem[16'h516B] = 8'h8D;
mem[16'h516C] = 8'hC0;
mem[16'h516D] = 8'h65;
mem[16'h516E] = 8'h20;
mem[16'h516F] = 8'h6A;
mem[16'h5170] = 8'h65;
mem[16'h5171] = 8'hA6;
mem[16'h5172] = 8'h70;
mem[16'h5173] = 8'hA9;
mem[16'h5174] = 8'h00;
mem[16'h5175] = 8'h9D;
mem[16'h5176] = 8'h1C;
mem[16'h5177] = 8'h51;
mem[16'h5178] = 8'h60;
mem[16'h5179] = 8'h01;
mem[16'h517A] = 8'h07;
mem[16'h517B] = 8'h1F;
mem[16'h517C] = 8'h1F;
mem[16'h517D] = 8'h1F;
mem[16'h517E] = 8'h1F;
mem[16'h517F] = 8'h1F;
mem[16'h5180] = 8'h07;
mem[16'h5181] = 8'h01;
mem[16'h5182] = 8'h1E;
mem[16'h5183] = 8'h00;
mem[16'h5184] = 8'h78;
mem[16'h5185] = 8'h00;
mem[16'h5186] = 8'h60;
mem[16'h5187] = 8'h03;
mem[16'h5188] = 8'h60;
mem[16'h5189] = 8'h03;
mem[16'h518A] = 8'h60;
mem[16'h518B] = 8'h03;
mem[16'h518C] = 8'h60;
mem[16'h518D] = 8'h03;
mem[16'h518E] = 8'h60;
mem[16'h518F] = 8'h03;
mem[16'h5190] = 8'h78;
mem[16'h5191] = 8'h00;
mem[16'h5192] = 8'h1E;
mem[16'h5193] = 8'h00;
mem[16'h5194] = 8'h06;
mem[16'h5195] = 8'h18;
mem[16'h5196] = 8'h60;
mem[16'h5197] = 8'h60;
mem[16'h5198] = 8'h60;
mem[16'h5199] = 8'h60;
mem[16'h519A] = 8'h60;
mem[16'h519B] = 8'h18;
mem[16'h519C] = 8'h06;
mem[16'h519D] = 8'hA9;
mem[16'h519E] = 8'h00;
mem[16'h519F] = 8'h8D;
mem[16'h51A0] = 8'h19;
mem[16'h51A1] = 8'h52;
mem[16'h51A2] = 8'h8D;
mem[16'h51A3] = 8'h8D;
mem[16'h51A4] = 8'h52;
mem[16'h51A5] = 8'h8D;
mem[16'h51A6] = 8'h8E;
mem[16'h51A7] = 8'h52;
mem[16'h51A8] = 8'h8D;
mem[16'h51A9] = 8'h8F;
mem[16'h51AA] = 8'h52;
mem[16'h51AB] = 8'h8D;
mem[16'h51AC] = 8'h90;
mem[16'h51AD] = 8'h52;
mem[16'h51AE] = 8'h8D;
mem[16'h51AF] = 8'h91;
mem[16'h51B0] = 8'h52;
mem[16'h51B1] = 8'h8D;
mem[16'h51B2] = 8'h92;
mem[16'h51B3] = 8'h52;
mem[16'h51B4] = 8'h8D;
mem[16'h51B5] = 8'h93;
mem[16'h51B6] = 8'h52;
mem[16'h51B7] = 8'h8D;
mem[16'h51B8] = 8'h94;
mem[16'h51B9] = 8'h52;
mem[16'h51BA] = 8'hA9;
mem[16'h51BB] = 8'h01;
mem[16'h51BC] = 8'h8D;
mem[16'h51BD] = 8'h1F;
mem[16'h51BE] = 8'h53;
mem[16'h51BF] = 8'h8D;
mem[16'h51C0] = 8'h20;
mem[16'h51C1] = 8'h53;
mem[16'h51C2] = 8'h8D;
mem[16'h51C3] = 8'h21;
mem[16'h51C4] = 8'h53;
mem[16'h51C5] = 8'h8D;
mem[16'h51C6] = 8'h22;
mem[16'h51C7] = 8'h53;
mem[16'h51C8] = 8'hAD;
mem[16'h51C9] = 8'h27;
mem[16'h51CA] = 8'h53;
mem[16'h51CB] = 8'h8D;
mem[16'h51CC] = 8'h28;
mem[16'h51CD] = 8'h53;
mem[16'h51CE] = 8'h8D;
mem[16'h51CF] = 8'h29;
mem[16'h51D0] = 8'h53;
mem[16'h51D1] = 8'h8D;
mem[16'h51D2] = 8'h2A;
mem[16'h51D3] = 8'h53;
mem[16'h51D4] = 8'h8D;
mem[16'h51D5] = 8'h2B;
mem[16'h51D6] = 8'h53;
mem[16'h51D7] = 8'hA9;
mem[16'h51D8] = 8'h01;
mem[16'h51D9] = 8'h8D;
mem[16'h51DA] = 8'h19;
mem[16'h51DB] = 8'h52;
mem[16'h51DC] = 8'h20;
mem[16'h51DD] = 8'h18;
mem[16'h51DE] = 8'h52;
mem[16'h51DF] = 8'hAD;
mem[16'h51E0] = 8'h1F;
mem[16'h51E1] = 8'h53;
mem[16'h51E2] = 8'hC9;
mem[16'h51E3] = 8'h4E;
mem[16'h51E4] = 8'h90;
mem[16'h51E5] = 8'hF6;
mem[16'h51E6] = 8'hA9;
mem[16'h51E7] = 8'h02;
mem[16'h51E8] = 8'h8D;
mem[16'h51E9] = 8'h19;
mem[16'h51EA] = 8'h52;
mem[16'h51EB] = 8'h20;
mem[16'h51EC] = 8'h18;
mem[16'h51ED] = 8'h52;
mem[16'h51EE] = 8'hAD;
mem[16'h51EF] = 8'h1F;
mem[16'h51F0] = 8'h53;
mem[16'h51F1] = 8'hC9;
mem[16'h51F2] = 8'hA4;
mem[16'h51F3] = 8'h90;
mem[16'h51F4] = 8'hF6;
mem[16'h51F5] = 8'hA9;
mem[16'h51F6] = 8'h03;
mem[16'h51F7] = 8'hCD;
mem[16'h51F8] = 8'hB3;
mem[16'h51F9] = 8'h4A;
mem[16'h51FA] = 8'hF0;
mem[16'h51FB] = 8'h02;
mem[16'h51FC] = 8'hB0;
mem[16'h51FD] = 8'h19;
mem[16'h51FE] = 8'h8D;
mem[16'h51FF] = 8'h19;
mem[16'h5200] = 8'h52;
mem[16'h5201] = 8'h20;
mem[16'h5202] = 8'h18;
mem[16'h5203] = 8'h52;
mem[16'h5204] = 8'hAD;
mem[16'h5205] = 8'h1F;
mem[16'h5206] = 8'h53;
mem[16'h5207] = 8'hC9;
mem[16'h5208] = 8'hF4;
mem[16'h5209] = 8'h90;
mem[16'h520A] = 8'hF6;
mem[16'h520B] = 8'hA9;
mem[16'h520C] = 8'h04;
mem[16'h520D] = 8'hCD;
mem[16'h520E] = 8'hB3;
mem[16'h520F] = 8'h4A;
mem[16'h5210] = 8'hF0;
mem[16'h5211] = 8'h02;
mem[16'h5212] = 8'hB0;
mem[16'h5213] = 8'h03;
mem[16'h5214] = 8'h8D;
mem[16'h5215] = 8'h19;
mem[16'h5216] = 8'h52;
mem[16'h5217] = 8'h60;
mem[16'h5218] = 8'hA2;
mem[16'h5219] = 8'h03;
mem[16'h521A] = 8'hCA;
mem[16'h521B] = 8'h30;
mem[16'h521C] = 8'h3F;
mem[16'h521D] = 8'h86;
mem[16'h521E] = 8'h70;
mem[16'h521F] = 8'h20;
mem[16'h5220] = 8'hEE;
mem[16'h5221] = 8'h52;
mem[16'h5222] = 8'hA6;
mem[16'h5223] = 8'h70;
mem[16'h5224] = 8'hBD;
mem[16'h5225] = 8'h1F;
mem[16'h5226] = 8'h53;
mem[16'h5227] = 8'hC9;
mem[16'h5228] = 8'hFD;
mem[16'h5229] = 8'hB0;
mem[16'h522A] = 8'h0E;
mem[16'h522B] = 8'h18;
mem[16'h522C] = 8'h69;
mem[16'h522D] = 8'h02;
mem[16'h522E] = 8'h9D;
mem[16'h522F] = 8'h1F;
mem[16'h5230] = 8'h53;
mem[16'h5231] = 8'h20;
mem[16'h5232] = 8'h5D;
mem[16'h5233] = 8'h52;
mem[16'h5234] = 8'hA6;
mem[16'h5235] = 8'h70;
mem[16'h5236] = 8'h4C;
mem[16'h5237] = 8'h1A;
mem[16'h5238] = 8'h52;
mem[16'h5239] = 8'hBD;
mem[16'h523A] = 8'h28;
mem[16'h523B] = 8'h53;
mem[16'h523C] = 8'h38;
mem[16'h523D] = 8'hE9;
mem[16'h523E] = 8'h02;
mem[16'h523F] = 8'h9D;
mem[16'h5240] = 8'h28;
mem[16'h5241] = 8'h53;
mem[16'h5242] = 8'hD0;
mem[16'h5243] = 8'hD6;
mem[16'h5244] = 8'h20;
mem[16'h5245] = 8'h64;
mem[16'h5246] = 8'h52;
mem[16'h5247] = 8'hA6;
mem[16'h5248] = 8'h70;
mem[16'h5249] = 8'hA9;
mem[16'h524A] = 8'h00;
mem[16'h524B] = 8'h9D;
mem[16'h524C] = 8'h8D;
mem[16'h524D] = 8'h52;
mem[16'h524E] = 8'hA9;
mem[16'h524F] = 8'h01;
mem[16'h5250] = 8'h9D;
mem[16'h5251] = 8'h1F;
mem[16'h5252] = 8'h53;
mem[16'h5253] = 8'hAD;
mem[16'h5254] = 8'h27;
mem[16'h5255] = 8'h53;
mem[16'h5256] = 8'h9D;
mem[16'h5257] = 8'h28;
mem[16'h5258] = 8'h53;
mem[16'h5259] = 8'h4C;
mem[16'h525A] = 8'h1A;
mem[16'h525B] = 8'h52;
mem[16'h525C] = 8'h60;
mem[16'h525D] = 8'hA6;
mem[16'h525E] = 8'h70;
mem[16'h525F] = 8'hBD;
mem[16'h5260] = 8'h8D;
mem[16'h5261] = 8'h52;
mem[16'h5262] = 8'hD0;
mem[16'h5263] = 8'h28;
mem[16'h5264] = 8'hA6;
mem[16'h5265] = 8'h70;
mem[16'h5266] = 8'hBD;
mem[16'h5267] = 8'h23;
mem[16'h5268] = 8'h53;
mem[16'h5269] = 8'h85;
mem[16'h526A] = 8'h56;
mem[16'h526B] = 8'hBD;
mem[16'h526C] = 8'h1F;
mem[16'h526D] = 8'h53;
mem[16'h526E] = 8'h38;
mem[16'h526F] = 8'hFD;
mem[16'h5270] = 8'h28;
mem[16'h5271] = 8'h53;
mem[16'h5272] = 8'h90;
mem[16'h5273] = 8'h18;
mem[16'h5274] = 8'h85;
mem[16'h5275] = 8'h57;
mem[16'h5276] = 8'hA9;
mem[16'h5277] = 8'h09;
mem[16'h5278] = 8'h8D;
mem[16'h5279] = 8'hC0;
mem[16'h527A] = 8'h65;
mem[16'h527B] = 8'hA9;
mem[16'h527C] = 8'hC9;
mem[16'h527D] = 8'hA0;
mem[16'h527E] = 8'h50;
mem[16'h527F] = 8'h20;
mem[16'h5280] = 8'hC7;
mem[16'h5281] = 8'h65;
mem[16'h5282] = 8'h20;
mem[16'h5283] = 8'h6A;
mem[16'h5284] = 8'h65;
mem[16'h5285] = 8'hA6;
mem[16'h5286] = 8'h70;
mem[16'h5287] = 8'hA9;
mem[16'h5288] = 8'h01;
mem[16'h5289] = 8'h9D;
mem[16'h528A] = 8'h8D;
mem[16'h528B] = 8'h52;
mem[16'h528C] = 8'h60;
mem[16'h528D] = 8'h01;
mem[16'h528E] = 8'h01;
mem[16'h528F] = 8'h01;
mem[16'h5290] = 8'h00;
mem[16'h5291] = 8'h09;
mem[16'h5292] = 8'h09;
mem[16'h5293] = 8'h09;
mem[16'h5294] = 8'h00;
mem[16'h5295] = 8'hBD;
mem[16'h5296] = 8'h91;
mem[16'h5297] = 8'h52;
mem[16'h5298] = 8'hD0;
mem[16'h5299] = 8'h12;
mem[16'h529A] = 8'hA9;
mem[16'h529B] = 8'h79;
mem[16'h529C] = 8'hA0;
mem[16'h529D] = 8'h51;
mem[16'h529E] = 8'h20;
mem[16'h529F] = 8'hC7;
mem[16'h52A0] = 8'h65;
mem[16'h52A1] = 8'hA9;
mem[16'h52A2] = 8'h09;
mem[16'h52A3] = 8'h8D;
mem[16'h52A4] = 8'hC0;
mem[16'h52A5] = 8'h65;
mem[16'h52A6] = 8'h9D;
mem[16'h52A7] = 8'h91;
mem[16'h52A8] = 8'h52;
mem[16'h52A9] = 8'h20;
mem[16'h52AA] = 8'h6A;
mem[16'h52AB] = 8'h65;
mem[16'h52AC] = 8'hA6;
mem[16'h52AD] = 8'h70;
mem[16'h52AE] = 8'hBD;
mem[16'h52AF] = 8'h23;
mem[16'h52B0] = 8'h53;
mem[16'h52B1] = 8'h85;
mem[16'h52B2] = 8'h56;
mem[16'h52B3] = 8'hBC;
mem[16'h52B4] = 8'h1F;
mem[16'h52B5] = 8'h53;
mem[16'h52B6] = 8'h84;
mem[16'h52B7] = 8'h57;
mem[16'h52B8] = 8'hB9;
mem[16'h52B9] = 8'h3E;
mem[16'h52BA] = 8'h8C;
mem[16'h52BB] = 8'hAA;
mem[16'h52BC] = 8'hBD;
mem[16'h52BD] = 8'h94;
mem[16'h52BE] = 8'h8E;
mem[16'h52BF] = 8'hAA;
mem[16'h52C0] = 8'hBD;
mem[16'h52C1] = 8'h66;
mem[16'h52C2] = 8'h62;
mem[16'h52C3] = 8'hBC;
mem[16'h52C4] = 8'h6D;
mem[16'h52C5] = 8'h62;
mem[16'h52C6] = 8'h20;
mem[16'h52C7] = 8'hF4;
mem[16'h52C8] = 8'h71;
mem[16'h52C9] = 8'hA9;
mem[16'h52CA] = 8'h12;
mem[16'h52CB] = 8'h8D;
mem[16'h52CC] = 8'hED;
mem[16'h52CD] = 8'h71;
mem[16'h52CE] = 8'h20;
mem[16'h52CF] = 8'hAC;
mem[16'h52D0] = 8'h71;
mem[16'h52D1] = 8'h60;
mem[16'h52D2] = 8'hBD;
mem[16'h52D3] = 8'h91;
mem[16'h52D4] = 8'h52;
mem[16'h52D5] = 8'hF0;
mem[16'h52D6] = 8'h16;
mem[16'h52D7] = 8'hA9;
mem[16'h52D8] = 8'h79;
mem[16'h52D9] = 8'hA0;
mem[16'h52DA] = 8'h51;
mem[16'h52DB] = 8'h20;
mem[16'h52DC] = 8'hC7;
mem[16'h52DD] = 8'h65;
mem[16'h52DE] = 8'hA9;
mem[16'h52DF] = 8'h09;
mem[16'h52E0] = 8'h8D;
mem[16'h52E1] = 8'hC0;
mem[16'h52E2] = 8'h65;
mem[16'h52E3] = 8'h20;
mem[16'h52E4] = 8'h6A;
mem[16'h52E5] = 8'h65;
mem[16'h52E6] = 8'hA6;
mem[16'h52E7] = 8'h70;
mem[16'h52E8] = 8'hA9;
mem[16'h52E9] = 8'h00;
mem[16'h52EA] = 8'h9D;
mem[16'h52EB] = 8'h91;
mem[16'h52EC] = 8'h52;
mem[16'h52ED] = 8'h60;
mem[16'h52EE] = 8'hA6;
mem[16'h52EF] = 8'h70;
mem[16'h52F0] = 8'hBD;
mem[16'h52F1] = 8'h23;
mem[16'h52F2] = 8'h53;
mem[16'h52F3] = 8'h85;
mem[16'h52F4] = 8'h56;
mem[16'h52F5] = 8'h85;
mem[16'h52F6] = 8'h6F;
mem[16'h52F7] = 8'hBD;
mem[16'h52F8] = 8'h1F;
mem[16'h52F9] = 8'h53;
mem[16'h52FA] = 8'h85;
mem[16'h52FB] = 8'h57;
mem[16'h52FC] = 8'hC9;
mem[16'h52FD] = 8'hFD;
mem[16'h52FE] = 8'hF0;
mem[16'h52FF] = 8'h08;
mem[16'h5300] = 8'hB0;
mem[16'h5301] = 8'h09;
mem[16'h5302] = 8'h20;
mem[16'h5303] = 8'h95;
mem[16'h5304] = 8'h52;
mem[16'h5305] = 8'h4C;
mem[16'h5306] = 8'h0B;
mem[16'h5307] = 8'h53;
mem[16'h5308] = 8'h20;
mem[16'h5309] = 8'hD2;
mem[16'h530A] = 8'h52;
mem[16'h530B] = 8'hA6;
mem[16'h530C] = 8'h70;
mem[16'h530D] = 8'hA5;
mem[16'h530E] = 8'h57;
mem[16'h530F] = 8'h38;
mem[16'h5310] = 8'hFD;
mem[16'h5311] = 8'h28;
mem[16'h5312] = 8'h53;
mem[16'h5313] = 8'h90;
mem[16'h5314] = 8'h09;
mem[16'h5315] = 8'h85;
mem[16'h5316] = 8'h57;
mem[16'h5317] = 8'hA5;
mem[16'h5318] = 8'h6F;
mem[16'h5319] = 8'h85;
mem[16'h531A] = 8'h56;
mem[16'h531B] = 8'h20;
mem[16'h531C] = 8'h99;
mem[16'h531D] = 8'h54;
mem[16'h531E] = 8'h60;
mem[16'h531F] = 8'hF5;
mem[16'h5320] = 8'hA7;
mem[16'h5321] = 8'h51;
mem[16'h5322] = 8'h01;
mem[16'h5323] = 8'h41;
mem[16'h5324] = 8'h41;
mem[16'h5325] = 8'h41;
mem[16'h5326] = 8'h41;
mem[16'h5327] = 8'h30;
mem[16'h5328] = 8'h30;
mem[16'h5329] = 8'h30;
mem[16'h532A] = 8'h30;
mem[16'h532B] = 8'h30;
mem[16'h532C] = 8'hAD;
mem[16'h532D] = 8'hB1;
mem[16'h532E] = 8'h4A;
mem[16'h532F] = 8'h8D;
mem[16'h5330] = 8'h8B;
mem[16'h5331] = 8'h53;
mem[16'h5332] = 8'hF0;
mem[16'h5333] = 8'h55;
mem[16'h5334] = 8'hA9;
mem[16'h5335] = 8'h00;
mem[16'h5336] = 8'h8D;
mem[16'h5337] = 8'h09;
mem[16'h5338] = 8'h54;
mem[16'h5339] = 8'h8D;
mem[16'h533A] = 8'h0A;
mem[16'h533B] = 8'h54;
mem[16'h533C] = 8'h8D;
mem[16'h533D] = 8'h0B;
mem[16'h533E] = 8'h54;
mem[16'h533F] = 8'h8D;
mem[16'h5340] = 8'h06;
mem[16'h5341] = 8'h54;
mem[16'h5342] = 8'h8D;
mem[16'h5343] = 8'h07;
mem[16'h5344] = 8'h54;
mem[16'h5345] = 8'h8D;
mem[16'h5346] = 8'h08;
mem[16'h5347] = 8'h54;
mem[16'h5348] = 8'hA9;
mem[16'h5349] = 8'h01;
mem[16'h534A] = 8'h8D;
mem[16'h534B] = 8'h00;
mem[16'h534C] = 8'h54;
mem[16'h534D] = 8'h8D;
mem[16'h534E] = 8'h01;
mem[16'h534F] = 8'h54;
mem[16'h5350] = 8'h8D;
mem[16'h5351] = 8'h02;
mem[16'h5352] = 8'h54;
mem[16'h5353] = 8'hAD;
mem[16'h5354] = 8'h0C;
mem[16'h5355] = 8'h54;
mem[16'h5356] = 8'h8D;
mem[16'h5357] = 8'h0D;
mem[16'h5358] = 8'h54;
mem[16'h5359] = 8'h8D;
mem[16'h535A] = 8'h0E;
mem[16'h535B] = 8'h54;
mem[16'h535C] = 8'h8D;
mem[16'h535D] = 8'h0F;
mem[16'h535E] = 8'h54;
mem[16'h535F] = 8'hA9;
mem[16'h5360] = 8'h01;
mem[16'h5361] = 8'h8D;
mem[16'h5362] = 8'h8B;
mem[16'h5363] = 8'h53;
mem[16'h5364] = 8'h20;
mem[16'h5365] = 8'h8A;
mem[16'h5366] = 8'h53;
mem[16'h5367] = 8'hAD;
mem[16'h5368] = 8'h00;
mem[16'h5369] = 8'h54;
mem[16'h536A] = 8'hC9;
mem[16'h536B] = 8'h56;
mem[16'h536C] = 8'h90;
mem[16'h536D] = 8'hF6;
mem[16'h536E] = 8'hA9;
mem[16'h536F] = 8'h02;
mem[16'h5370] = 8'h8D;
mem[16'h5371] = 8'h8B;
mem[16'h5372] = 8'h53;
mem[16'h5373] = 8'h20;
mem[16'h5374] = 8'h8A;
mem[16'h5375] = 8'h53;
mem[16'h5376] = 8'hAD;
mem[16'h5377] = 8'h00;
mem[16'h5378] = 8'h54;
mem[16'h5379] = 8'hC9;
mem[16'h537A] = 8'hC0;
mem[16'h537B] = 8'h90;
mem[16'h537C] = 8'hF6;
mem[16'h537D] = 8'hA9;
mem[16'h537E] = 8'h03;
mem[16'h537F] = 8'hCD;
mem[16'h5380] = 8'hB1;
mem[16'h5381] = 8'h4A;
mem[16'h5382] = 8'hF0;
mem[16'h5383] = 8'h02;
mem[16'h5384] = 8'hB0;
mem[16'h5385] = 8'h03;
mem[16'h5386] = 8'h8D;
mem[16'h5387] = 8'h8B;
mem[16'h5388] = 8'h53;
mem[16'h5389] = 8'h60;
mem[16'h538A] = 8'hA2;
mem[16'h538B] = 8'h03;
mem[16'h538C] = 8'hCA;
mem[16'h538D] = 8'h30;
mem[16'h538E] = 8'h3F;
mem[16'h538F] = 8'h86;
mem[16'h5390] = 8'h70;
mem[16'h5391] = 8'h20;
mem[16'h5392] = 8'hCF;
mem[16'h5393] = 8'h53;
mem[16'h5394] = 8'hA6;
mem[16'h5395] = 8'h70;
mem[16'h5396] = 8'hBD;
mem[16'h5397] = 8'h00;
mem[16'h5398] = 8'h54;
mem[16'h5399] = 8'hC9;
mem[16'h539A] = 8'hFD;
mem[16'h539B] = 8'hB0;
mem[16'h539C] = 8'h0E;
mem[16'h539D] = 8'h18;
mem[16'h539E] = 8'h69;
mem[16'h539F] = 8'h02;
mem[16'h53A0] = 8'h9D;
mem[16'h53A1] = 8'h00;
mem[16'h53A2] = 8'h54;
mem[16'h53A3] = 8'h20;
mem[16'h53A4] = 8'h69;
mem[16'h53A5] = 8'h54;
mem[16'h53A6] = 8'hA6;
mem[16'h53A7] = 8'h70;
mem[16'h53A8] = 8'h4C;
mem[16'h53A9] = 8'h8C;
mem[16'h53AA] = 8'h53;
mem[16'h53AB] = 8'hBD;
mem[16'h53AC] = 8'h0D;
mem[16'h53AD] = 8'h54;
mem[16'h53AE] = 8'h38;
mem[16'h53AF] = 8'hE9;
mem[16'h53B0] = 8'h02;
mem[16'h53B1] = 8'h9D;
mem[16'h53B2] = 8'h0D;
mem[16'h53B3] = 8'h54;
mem[16'h53B4] = 8'hD0;
mem[16'h53B5] = 8'hD6;
mem[16'h53B6] = 8'h20;
mem[16'h53B7] = 8'h70;
mem[16'h53B8] = 8'h54;
mem[16'h53B9] = 8'hA6;
mem[16'h53BA] = 8'h70;
mem[16'h53BB] = 8'hA9;
mem[16'h53BC] = 8'h00;
mem[16'h53BD] = 8'h9D;
mem[16'h53BE] = 8'h09;
mem[16'h53BF] = 8'h54;
mem[16'h53C0] = 8'hA9;
mem[16'h53C1] = 8'h01;
mem[16'h53C2] = 8'h9D;
mem[16'h53C3] = 8'h00;
mem[16'h53C4] = 8'h54;
mem[16'h53C5] = 8'hAD;
mem[16'h53C6] = 8'h0C;
mem[16'h53C7] = 8'h54;
mem[16'h53C8] = 8'h9D;
mem[16'h53C9] = 8'h0D;
mem[16'h53CA] = 8'h54;
mem[16'h53CB] = 8'h4C;
mem[16'h53CC] = 8'h8C;
mem[16'h53CD] = 8'h53;
mem[16'h53CE] = 8'h60;
mem[16'h53CF] = 8'hA6;
mem[16'h53D0] = 8'h70;
mem[16'h53D1] = 8'hBD;
mem[16'h53D2] = 8'h03;
mem[16'h53D3] = 8'h54;
mem[16'h53D4] = 8'h85;
mem[16'h53D5] = 8'h56;
mem[16'h53D6] = 8'h85;
mem[16'h53D7] = 8'h6F;
mem[16'h53D8] = 8'hBD;
mem[16'h53D9] = 8'h00;
mem[16'h53DA] = 8'h54;
mem[16'h53DB] = 8'h85;
mem[16'h53DC] = 8'h57;
mem[16'h53DD] = 8'hC9;
mem[16'h53DE] = 8'hFD;
mem[16'h53DF] = 8'hF0;
mem[16'h53E0] = 8'h08;
mem[16'h53E1] = 8'hB0;
mem[16'h53E2] = 8'h09;
mem[16'h53E3] = 8'h20;
mem[16'h53E4] = 8'h10;
mem[16'h53E5] = 8'h54;
mem[16'h53E6] = 8'h4C;
mem[16'h53E7] = 8'hEC;
mem[16'h53E8] = 8'h53;
mem[16'h53E9] = 8'h20;
mem[16'h53EA] = 8'h4D;
mem[16'h53EB] = 8'h54;
mem[16'h53EC] = 8'hA6;
mem[16'h53ED] = 8'h70;
mem[16'h53EE] = 8'hA5;
mem[16'h53EF] = 8'h57;
mem[16'h53F0] = 8'h38;
mem[16'h53F1] = 8'hFD;
mem[16'h53F2] = 8'h0D;
mem[16'h53F3] = 8'h54;
mem[16'h53F4] = 8'h90;
mem[16'h53F5] = 8'h09;
mem[16'h53F6] = 8'h85;
mem[16'h53F7] = 8'h57;
mem[16'h53F8] = 8'hA5;
mem[16'h53F9] = 8'h6F;
mem[16'h53FA] = 8'h85;
mem[16'h53FB] = 8'h56;
mem[16'h53FC] = 8'h20;
mem[16'h53FD] = 8'h99;
mem[16'h53FE] = 8'h54;
mem[16'h53FF] = 8'h60;
mem[16'h5400] = 8'hC1;
mem[16'h5401] = 8'h6B;
mem[16'h5402] = 8'h01;
mem[16'h5403] = 8'h17;
mem[16'h5404] = 8'h17;
mem[16'h5405] = 8'h17;
mem[16'h5406] = 8'h09;
mem[16'h5407] = 8'h09;
mem[16'h5408] = 8'h00;
mem[16'h5409] = 8'h01;
mem[16'h540A] = 8'h01;
mem[16'h540B] = 8'h00;
mem[16'h540C] = 8'h40;
mem[16'h540D] = 8'h40;
mem[16'h540E] = 8'h40;
mem[16'h540F] = 8'h40;
mem[16'h5410] = 8'hBD;
mem[16'h5411] = 8'h06;
mem[16'h5412] = 8'h54;
mem[16'h5413] = 8'hD0;
mem[16'h5414] = 8'h12;
mem[16'h5415] = 8'hA9;
mem[16'h5416] = 8'h79;
mem[16'h5417] = 8'hA0;
mem[16'h5418] = 8'h51;
mem[16'h5419] = 8'h20;
mem[16'h541A] = 8'hC7;
mem[16'h541B] = 8'h65;
mem[16'h541C] = 8'hA9;
mem[16'h541D] = 8'h09;
mem[16'h541E] = 8'h8D;
mem[16'h541F] = 8'hC0;
mem[16'h5420] = 8'h65;
mem[16'h5421] = 8'h9D;
mem[16'h5422] = 8'h06;
mem[16'h5423] = 8'h54;
mem[16'h5424] = 8'h20;
mem[16'h5425] = 8'h6A;
mem[16'h5426] = 8'h65;
mem[16'h5427] = 8'hA6;
mem[16'h5428] = 8'h70;
mem[16'h5429] = 8'hBD;
mem[16'h542A] = 8'h03;
mem[16'h542B] = 8'h54;
mem[16'h542C] = 8'h85;
mem[16'h542D] = 8'h56;
mem[16'h542E] = 8'hBC;
mem[16'h542F] = 8'h00;
mem[16'h5430] = 8'h54;
mem[16'h5431] = 8'h84;
mem[16'h5432] = 8'h57;
mem[16'h5433] = 8'hB9;
mem[16'h5434] = 8'h3E;
mem[16'h5435] = 8'h8C;
mem[16'h5436] = 8'hAA;
mem[16'h5437] = 8'hBD;
mem[16'h5438] = 8'h94;
mem[16'h5439] = 8'h8E;
mem[16'h543A] = 8'hAA;
mem[16'h543B] = 8'hBD;
mem[16'h543C] = 8'h66;
mem[16'h543D] = 8'h62;
mem[16'h543E] = 8'hBC;
mem[16'h543F] = 8'h6D;
mem[16'h5440] = 8'h62;
mem[16'h5441] = 8'h20;
mem[16'h5442] = 8'hF4;
mem[16'h5443] = 8'h71;
mem[16'h5444] = 8'hA9;
mem[16'h5445] = 8'h12;
mem[16'h5446] = 8'h8D;
mem[16'h5447] = 8'hED;
mem[16'h5448] = 8'h71;
mem[16'h5449] = 8'h20;
mem[16'h544A] = 8'hAC;
mem[16'h544B] = 8'h71;
mem[16'h544C] = 8'h60;
mem[16'h544D] = 8'hBD;
mem[16'h544E] = 8'h06;
mem[16'h544F] = 8'h54;
mem[16'h5450] = 8'hF0;
mem[16'h5451] = 8'h16;
mem[16'h5452] = 8'hA9;
mem[16'h5453] = 8'h79;
mem[16'h5454] = 8'hA0;
mem[16'h5455] = 8'h51;
mem[16'h5456] = 8'h20;
mem[16'h5457] = 8'hC7;
mem[16'h5458] = 8'h65;
mem[16'h5459] = 8'hA9;
mem[16'h545A] = 8'h09;
mem[16'h545B] = 8'h8D;
mem[16'h545C] = 8'hC0;
mem[16'h545D] = 8'h65;
mem[16'h545E] = 8'h20;
mem[16'h545F] = 8'h6A;
mem[16'h5460] = 8'h65;
mem[16'h5461] = 8'hA6;
mem[16'h5462] = 8'h70;
mem[16'h5463] = 8'hA9;
mem[16'h5464] = 8'h00;
mem[16'h5465] = 8'h9D;
mem[16'h5466] = 8'h06;
mem[16'h5467] = 8'h54;
mem[16'h5468] = 8'h60;
mem[16'h5469] = 8'hA6;
mem[16'h546A] = 8'h70;
mem[16'h546B] = 8'hBD;
mem[16'h546C] = 8'h09;
mem[16'h546D] = 8'h54;
mem[16'h546E] = 8'hD0;
mem[16'h546F] = 8'h28;
mem[16'h5470] = 8'hA6;
mem[16'h5471] = 8'h70;
mem[16'h5472] = 8'hBD;
mem[16'h5473] = 8'h03;
mem[16'h5474] = 8'h54;
mem[16'h5475] = 8'h85;
mem[16'h5476] = 8'h56;
mem[16'h5477] = 8'hBD;
mem[16'h5478] = 8'h00;
mem[16'h5479] = 8'h54;
mem[16'h547A] = 8'h38;
mem[16'h547B] = 8'hFD;
mem[16'h547C] = 8'h0D;
mem[16'h547D] = 8'h54;
mem[16'h547E] = 8'h90;
mem[16'h547F] = 8'h18;
mem[16'h5480] = 8'h85;
mem[16'h5481] = 8'h57;
mem[16'h5482] = 8'hA9;
mem[16'h5483] = 8'h09;
mem[16'h5484] = 8'h8D;
mem[16'h5485] = 8'hC0;
mem[16'h5486] = 8'h65;
mem[16'h5487] = 8'hA9;
mem[16'h5488] = 8'hC9;
mem[16'h5489] = 8'hA0;
mem[16'h548A] = 8'h50;
mem[16'h548B] = 8'h20;
mem[16'h548C] = 8'hC7;
mem[16'h548D] = 8'h65;
mem[16'h548E] = 8'h20;
mem[16'h548F] = 8'h6A;
mem[16'h5490] = 8'h65;
mem[16'h5491] = 8'hA9;
mem[16'h5492] = 8'h01;
mem[16'h5493] = 8'hA6;
mem[16'h5494] = 8'h70;
mem[16'h5495] = 8'h9D;
mem[16'h5496] = 8'h09;
mem[16'h5497] = 8'h54;
mem[16'h5498] = 8'h60;
mem[16'h5499] = 8'hA9;
mem[16'h549A] = 8'h09;
mem[16'h549B] = 8'h8D;
mem[16'h549C] = 8'hC0;
mem[16'h549D] = 8'h65;
mem[16'h549E] = 8'hA9;
mem[16'h549F] = 8'hA9;
mem[16'h54A0] = 8'hA0;
mem[16'h54A1] = 8'h54;
mem[16'h54A2] = 8'h20;
mem[16'h54A3] = 8'hC7;
mem[16'h54A4] = 8'h65;
mem[16'h54A5] = 8'h20;
mem[16'h54A6] = 8'h6A;
mem[16'h54A7] = 8'h65;
mem[16'h54A8] = 8'h60;
mem[16'h54A9] = 8'h30;
mem[16'h54AA] = 8'h0C;
mem[16'h54AB] = 8'h03;
mem[16'h54AC] = 8'h03;
mem[16'h54AD] = 8'h03;
mem[16'h54AE] = 8'h03;
mem[16'h54AF] = 8'h03;
mem[16'h54B0] = 8'h0C;
mem[16'h54B1] = 8'h30;
mem[16'h54B2] = 8'h85;
mem[16'h54B3] = 8'h57;
mem[16'h54B4] = 8'hA9;
mem[16'h54B5] = 8'h09;
mem[16'h54B6] = 8'h85;
mem[16'h54B7] = 8'h56;
mem[16'h54B8] = 8'hA4;
mem[16'h54B9] = 8'h56;
mem[16'h54BA] = 8'hB9;
mem[16'h54BB] = 8'hD5;
mem[16'h54BC] = 8'h8E;
mem[16'h54BD] = 8'h85;
mem[16'h54BE] = 8'h59;
mem[16'h54BF] = 8'hB9;
mem[16'h54C0] = 8'h95;
mem[16'h54C1] = 8'h8F;
mem[16'h54C2] = 8'h85;
mem[16'h54C3] = 8'h5A;
mem[16'h54C4] = 8'hA6;
mem[16'h54C5] = 8'h57;
mem[16'h54C6] = 8'hBC;
mem[16'h54C7] = 8'h56;
mem[16'h54C8] = 8'h8D;
mem[16'h54C9] = 8'hA5;
mem[16'h54CA] = 8'h57;
mem[16'h54CB] = 8'h29;
mem[16'h54CC] = 8'h01;
mem[16'h54CD] = 8'hF0;
mem[16'h54CE] = 8'h0D;
mem[16'h54CF] = 8'hA9;
mem[16'h54D0] = 8'hAA;
mem[16'h54D1] = 8'h8D;
mem[16'h54D2] = 8'hFA;
mem[16'h54D3] = 8'h54;
mem[16'h54D4] = 8'hA9;
mem[16'h54D5] = 8'hD5;
mem[16'h54D6] = 8'h8D;
mem[16'h54D7] = 8'hFB;
mem[16'h54D8] = 8'h54;
mem[16'h54D9] = 8'h4C;
mem[16'h54DA] = 8'hE6;
mem[16'h54DB] = 8'h54;
mem[16'h54DC] = 8'hA9;
mem[16'h54DD] = 8'hD5;
mem[16'h54DE] = 8'h8D;
mem[16'h54DF] = 8'hFA;
mem[16'h54E0] = 8'h54;
mem[16'h54E1] = 8'hA9;
mem[16'h54E2] = 8'hAA;
mem[16'h54E3] = 8'h8D;
mem[16'h54E4] = 8'hFB;
mem[16'h54E5] = 8'h54;
mem[16'h54E6] = 8'hAD;
mem[16'h54E7] = 8'hFA;
mem[16'h54E8] = 8'h54;
mem[16'h54E9] = 8'h91;
mem[16'h54EA] = 8'h59;
mem[16'h54EB] = 8'hC8;
mem[16'h54EC] = 8'hAD;
mem[16'h54ED] = 8'hFB;
mem[16'h54EE] = 8'h54;
mem[16'h54EF] = 8'h91;
mem[16'h54F0] = 8'h59;
mem[16'h54F1] = 8'hE6;
mem[16'h54F2] = 8'h56;
mem[16'h54F3] = 8'hA5;
mem[16'h54F4] = 8'h56;
mem[16'h54F5] = 8'hC9;
mem[16'h54F6] = 8'h15;
mem[16'h54F7] = 8'h90;
mem[16'h54F8] = 8'hBF;
mem[16'h54F9] = 8'h60;
mem[16'h54FA] = 8'hAA;
mem[16'h54FB] = 8'hD5;
mem[16'h54FC] = 8'hA9;
mem[16'h54FD] = 8'h16;
mem[16'h54FE] = 8'hA0;
mem[16'h54FF] = 8'h55;
mem[16'h5500] = 8'h20;
mem[16'h5501] = 8'hC7;
mem[16'h5502] = 8'h65;
mem[16'h5503] = 8'hAD;
mem[16'h5504] = 8'hA1;
mem[16'h5505] = 8'h55;
mem[16'h5506] = 8'h85;
mem[16'h5507] = 8'h57;
mem[16'h5508] = 8'hAD;
mem[16'h5509] = 8'hA2;
mem[16'h550A] = 8'h55;
mem[16'h550B] = 8'h85;
mem[16'h550C] = 8'h56;
mem[16'h550D] = 8'hA9;
mem[16'h550E] = 8'h05;
mem[16'h550F] = 8'h8D;
mem[16'h5510] = 8'hC0;
mem[16'h5511] = 8'h65;
mem[16'h5512] = 8'h20;
mem[16'h5513] = 8'h6A;
mem[16'h5514] = 8'h65;
mem[16'h5515] = 8'h60;
mem[16'h5516] = 8'hD5;
mem[16'h5517] = 8'hD5;
mem[16'h5518] = 8'hD5;
mem[16'h5519] = 8'hD5;
mem[16'h551A] = 8'hD5;
mem[16'h551B] = 8'hD5;
mem[16'h551C] = 8'hAA;
mem[16'h551D] = 8'hD5;
mem[16'h551E] = 8'hAA;
mem[16'h551F] = 8'hD5;
mem[16'h5520] = 8'hAA;
mem[16'h5521] = 8'hD5;
mem[16'h5522] = 8'hAA;
mem[16'h5523] = 8'hD5;
mem[16'h5524] = 8'hAA;
mem[16'h5525] = 8'hA9;
mem[16'h5526] = 8'h14;
mem[16'h5527] = 8'h8D;
mem[16'h5528] = 8'hA2;
mem[16'h5529] = 8'h55;
mem[16'h552A] = 8'hA9;
mem[16'h552B] = 8'h00;
mem[16'h552C] = 8'h8D;
mem[16'h552D] = 8'hA1;
mem[16'h552E] = 8'h55;
mem[16'h552F] = 8'h20;
mem[16'h5530] = 8'hFC;
mem[16'h5531] = 8'h54;
mem[16'h5532] = 8'hAD;
mem[16'h5533] = 8'hA1;
mem[16'h5534] = 8'h55;
mem[16'h5535] = 8'h18;
mem[16'h5536] = 8'h69;
mem[16'h5537] = 8'h08;
mem[16'h5538] = 8'hB0;
mem[16'h5539] = 8'h06;
mem[16'h553A] = 8'h8D;
mem[16'h553B] = 8'hA1;
mem[16'h553C] = 8'h55;
mem[16'h553D] = 8'h4C;
mem[16'h553E] = 8'h2F;
mem[16'h553F] = 8'h55;
mem[16'h5540] = 8'hAD;
mem[16'h5541] = 8'hA2;
mem[16'h5542] = 8'h55;
mem[16'h5543] = 8'h18;
mem[16'h5544] = 8'h69;
mem[16'h5545] = 8'h05;
mem[16'h5546] = 8'hC9;
mem[16'h5547] = 8'h56;
mem[16'h5548] = 8'hB0;
mem[16'h5549] = 8'h06;
mem[16'h554A] = 8'h8D;
mem[16'h554B] = 8'hA2;
mem[16'h554C] = 8'h55;
mem[16'h554D] = 8'h4C;
mem[16'h554E] = 8'h2A;
mem[16'h554F] = 8'h55;
mem[16'h5550] = 8'h60;
mem[16'h5551] = 8'hA9;
mem[16'h5552] = 8'h9B;
mem[16'h5553] = 8'hA0;
mem[16'h5554] = 8'h55;
mem[16'h5555] = 8'h20;
mem[16'h5556] = 8'hC7;
mem[16'h5557] = 8'h65;
mem[16'h5558] = 8'hA0;
mem[16'h5559] = 8'h04;
mem[16'h555A] = 8'hAE;
mem[16'h555B] = 8'hA0;
mem[16'h555C] = 8'h55;
mem[16'h555D] = 8'hB9;
mem[16'h555E] = 8'h8F;
mem[16'h555F] = 8'h55;
mem[16'h5560] = 8'h3D;
mem[16'h5561] = 8'h94;
mem[16'h5562] = 8'h55;
mem[16'h5563] = 8'h99;
mem[16'h5564] = 8'h9B;
mem[16'h5565] = 8'h55;
mem[16'h5566] = 8'hCE;
mem[16'h5567] = 8'hA0;
mem[16'h5568] = 8'h55;
mem[16'h5569] = 8'h10;
mem[16'h556A] = 8'h05;
mem[16'h556B] = 8'hA9;
mem[16'h556C] = 8'h06;
mem[16'h556D] = 8'h8D;
mem[16'h556E] = 8'hA0;
mem[16'h556F] = 8'h55;
mem[16'h5570] = 8'h88;
mem[16'h5571] = 8'h10;
mem[16'h5572] = 8'hE7;
mem[16'h5573] = 8'hA9;
mem[16'h5574] = 8'h05;
mem[16'h5575] = 8'h8D;
mem[16'h5576] = 8'hC0;
mem[16'h5577] = 8'h65;
mem[16'h5578] = 8'hAD;
mem[16'h5579] = 8'hA1;
mem[16'h557A] = 8'h55;
mem[16'h557B] = 8'h85;
mem[16'h557C] = 8'h57;
mem[16'h557D] = 8'hAD;
mem[16'h557E] = 8'hA2;
mem[16'h557F] = 8'h55;
mem[16'h5580] = 8'h85;
mem[16'h5581] = 8'h56;
mem[16'h5582] = 8'hC9;
mem[16'h5583] = 8'h12;
mem[16'h5584] = 8'hD0;
mem[16'h5585] = 8'h05;
mem[16'h5586] = 8'hA9;
mem[16'h5587] = 8'h02;
mem[16'h5588] = 8'h8D;
mem[16'h5589] = 8'hC0;
mem[16'h558A] = 8'h65;
mem[16'h558B] = 8'h20;
mem[16'h558C] = 8'h6A;
mem[16'h558D] = 8'h65;
mem[16'h558E] = 8'h60;
mem[16'h558F] = 8'h55;
mem[16'h5590] = 8'h55;
mem[16'h5591] = 8'h55;
mem[16'h5592] = 8'h55;
mem[16'h5593] = 8'h55;
mem[16'h5594] = 8'h51;
mem[16'h5595] = 8'h41;
mem[16'h5596] = 8'h45;
mem[16'h5597] = 8'h15;
mem[16'h5598] = 8'h54;
mem[16'h5599] = 8'h55;
mem[16'h559A] = 8'h05;
mem[16'h559B] = 8'h45;
mem[16'h559C] = 8'h15;
mem[16'h559D] = 8'h54;
mem[16'h559E] = 8'h55;
mem[16'h559F] = 8'h05;
mem[16'h55A0] = 8'h01;
mem[16'h55A1] = 8'h01;
mem[16'h55A2] = 8'h12;
mem[16'h55A3] = 8'hA9;
mem[16'h55A4] = 8'hAF;
mem[16'h55A5] = 8'h8D;
mem[16'h55A6] = 8'hA2;
mem[16'h55A7] = 8'h55;
mem[16'h55A8] = 8'hA9;
mem[16'h55A9] = 8'h00;
mem[16'h55AA] = 8'h8D;
mem[16'h55AB] = 8'hD8;
mem[16'h55AC] = 8'h77;
mem[16'h55AD] = 8'hA9;
mem[16'h55AE] = 8'h01;
mem[16'h55AF] = 8'h8D;
mem[16'h55B0] = 8'hA1;
mem[16'h55B1] = 8'h55;
mem[16'h55B2] = 8'h20;
mem[16'h55B3] = 8'h51;
mem[16'h55B4] = 8'h55;
mem[16'h55B5] = 8'hAD;
mem[16'h55B6] = 8'hA1;
mem[16'h55B7] = 8'h55;
mem[16'h55B8] = 8'h18;
mem[16'h55B9] = 8'h69;
mem[16'h55BA] = 8'h08;
mem[16'h55BB] = 8'hB0;
mem[16'h55BC] = 8'h06;
mem[16'h55BD] = 8'h8D;
mem[16'h55BE] = 8'hA1;
mem[16'h55BF] = 8'h55;
mem[16'h55C0] = 8'h4C;
mem[16'h55C1] = 8'hB2;
mem[16'h55C2] = 8'h55;
mem[16'h55C3] = 8'hAD;
mem[16'h55C4] = 8'hA2;
mem[16'h55C5] = 8'h55;
mem[16'h55C6] = 8'h18;
mem[16'h55C7] = 8'h69;
mem[16'h55C8] = 8'h05;
mem[16'h55C9] = 8'hC9;
mem[16'h55CA] = 8'hBE;
mem[16'h55CB] = 8'hB0;
mem[16'h55CC] = 8'h06;
mem[16'h55CD] = 8'h8D;
mem[16'h55CE] = 8'hA2;
mem[16'h55CF] = 8'h55;
mem[16'h55D0] = 8'h4C;
mem[16'h55D1] = 8'hAD;
mem[16'h55D2] = 8'h55;
mem[16'h55D3] = 8'hA9;
mem[16'h55D4] = 8'h5A;
mem[16'h55D5] = 8'h8D;
mem[16'h55D6] = 8'hA2;
mem[16'h55D7] = 8'h55;
mem[16'h55D8] = 8'hA9;
mem[16'h55D9] = 8'h01;
mem[16'h55DA] = 8'h8D;
mem[16'h55DB] = 8'hA1;
mem[16'h55DC] = 8'h55;
mem[16'h55DD] = 8'h20;
mem[16'h55DE] = 8'h51;
mem[16'h55DF] = 8'h55;
mem[16'h55E0] = 8'hAD;
mem[16'h55E1] = 8'hA1;
mem[16'h55E2] = 8'h55;
mem[16'h55E3] = 8'h18;
mem[16'h55E4] = 8'h69;
mem[16'h55E5] = 8'h08;
mem[16'h55E6] = 8'hB0;
mem[16'h55E7] = 8'h06;
mem[16'h55E8] = 8'h8D;
mem[16'h55E9] = 8'hA1;
mem[16'h55EA] = 8'h55;
mem[16'h55EB] = 8'h4C;
mem[16'h55EC] = 8'hDD;
mem[16'h55ED] = 8'h55;
mem[16'h55EE] = 8'hAD;
mem[16'h55EF] = 8'hA2;
mem[16'h55F0] = 8'h55;
mem[16'h55F1] = 8'h18;
mem[16'h55F2] = 8'h69;
mem[16'h55F3] = 8'h05;
mem[16'h55F4] = 8'hC9;
mem[16'h55F5] = 8'h65;
mem[16'h55F6] = 8'hB0;
mem[16'h55F7] = 8'h06;
mem[16'h55F8] = 8'h8D;
mem[16'h55F9] = 8'hA2;
mem[16'h55FA] = 8'h55;
mem[16'h55FB] = 8'h4C;
mem[16'h55FC] = 8'hD8;
mem[16'h55FD] = 8'h55;
mem[16'h55FE] = 8'h60;
mem[16'h55FF] = 8'hAE;
mem[16'h5600] = 8'hAE;
mem[16'h5601] = 8'h4A;
mem[16'h5602] = 8'hCA;
mem[16'h5603] = 8'h30;
mem[16'h5604] = 8'h29;
mem[16'h5605] = 8'h86;
mem[16'h5606] = 8'h70;
mem[16'h5607] = 8'hBD;
mem[16'h5608] = 8'h47;
mem[16'h5609] = 8'h60;
mem[16'h560A] = 8'hC9;
mem[16'h560B] = 8'h02;
mem[16'h560C] = 8'h90;
mem[16'h560D] = 8'h0E;
mem[16'h560E] = 8'h38;
mem[16'h560F] = 8'hE9;
mem[16'h5610] = 8'h02;
mem[16'h5611] = 8'h9D;
mem[16'h5612] = 8'h47;
mem[16'h5613] = 8'h60;
mem[16'h5614] = 8'h20;
mem[16'h5615] = 8'h2F;
mem[16'h5616] = 8'h56;
mem[16'h5617] = 8'hA6;
mem[16'h5618] = 8'h70;
mem[16'h5619] = 8'h4C;
mem[16'h561A] = 8'h02;
mem[16'h561B] = 8'h56;
mem[16'h561C] = 8'h20;
mem[16'h561D] = 8'h13;
mem[16'h561E] = 8'h60;
mem[16'h561F] = 8'hA6;
mem[16'h5620] = 8'h70;
mem[16'h5621] = 8'hA9;
mem[16'h5622] = 8'hFE;
mem[16'h5623] = 8'h9D;
mem[16'h5624] = 8'h47;
mem[16'h5625] = 8'h60;
mem[16'h5626] = 8'h20;
mem[16'h5627] = 8'h13;
mem[16'h5628] = 8'h60;
mem[16'h5629] = 8'hA6;
mem[16'h562A] = 8'h70;
mem[16'h562B] = 8'h4C;
mem[16'h562C] = 8'h02;
mem[16'h562D] = 8'h56;
mem[16'h562E] = 8'h60;
mem[16'h562F] = 8'hA6;
mem[16'h5630] = 8'h70;
mem[16'h5631] = 8'hBD;
mem[16'h5632] = 8'h4A;
mem[16'h5633] = 8'h60;
mem[16'h5634] = 8'h85;
mem[16'h5635] = 8'h56;
mem[16'h5636] = 8'hBC;
mem[16'h5637] = 8'h47;
mem[16'h5638] = 8'h60;
mem[16'h5639] = 8'h84;
mem[16'h563A] = 8'h57;
mem[16'h563B] = 8'hB9;
mem[16'h563C] = 8'h3E;
mem[16'h563D] = 8'h8C;
mem[16'h563E] = 8'hAA;
mem[16'h563F] = 8'hBD;
mem[16'h5640] = 8'h94;
mem[16'h5641] = 8'h8E;
mem[16'h5642] = 8'hAA;
mem[16'h5643] = 8'hBD;
mem[16'h5644] = 8'h55;
mem[16'h5645] = 8'h56;
mem[16'h5646] = 8'hBC;
mem[16'h5647] = 8'h5C;
mem[16'h5648] = 8'h56;
mem[16'h5649] = 8'h20;
mem[16'h564A] = 8'hD1;
mem[16'h564B] = 8'h8A;
mem[16'h564C] = 8'hA9;
mem[16'h564D] = 8'h20;
mem[16'h564E] = 8'h8D;
mem[16'h564F] = 8'hCA;
mem[16'h5650] = 8'h8A;
mem[16'h5651] = 8'h20;
mem[16'h5652] = 8'h79;
mem[16'h5653] = 8'h8A;
mem[16'h5654] = 8'h60;
mem[16'h5655] = 8'h63;
mem[16'h5656] = 8'h83;
mem[16'h5657] = 8'hA3;
mem[16'h5658] = 8'hC3;
mem[16'h5659] = 8'hE3;
mem[16'h565A] = 8'h03;
mem[16'h565B] = 8'h23;
mem[16'h565C] = 8'h56;
mem[16'h565D] = 8'h56;
mem[16'h565E] = 8'h56;
mem[16'h565F] = 8'h56;
mem[16'h5660] = 8'h56;
mem[16'h5661] = 8'h57;
mem[16'h5662] = 8'h57;
mem[16'h5663] = 8'h00;
mem[16'h5664] = 8'h0F;
mem[16'h5665] = 8'h3C;
mem[16'h5666] = 8'h00;
mem[16'h5667] = 8'h66;
mem[16'h5668] = 8'h01;
mem[16'h5669] = 8'h20;
mem[16'h566A] = 8'h00;
mem[16'h566B] = 8'h69;
mem[16'h566C] = 8'h01;
mem[16'h566D] = 8'h20;
mem[16'h566E] = 8'h00;
mem[16'h566F] = 8'h09;
mem[16'h5670] = 8'h02;
mem[16'h5671] = 8'h20;
mem[16'h5672] = 8'h00;
mem[16'h5673] = 8'h09;
mem[16'h5674] = 8'h02;
mem[16'h5675] = 8'h20;
mem[16'h5676] = 8'h00;
mem[16'h5677] = 8'h69;
mem[16'h5678] = 8'h01;
mem[16'h5679] = 8'h20;
mem[16'h567A] = 8'h00;
mem[16'h567B] = 8'h66;
mem[16'h567C] = 8'h01;
mem[16'h567D] = 8'h20;
mem[16'h567E] = 8'h00;
mem[16'h567F] = 8'h00;
mem[16'h5680] = 8'h0F;
mem[16'h5681] = 8'h3C;
mem[16'h5682] = 8'h00;
mem[16'h5683] = 8'h00;
mem[16'h5684] = 8'h1E;
mem[16'h5685] = 8'h78;
mem[16'h5686] = 8'h00;
mem[16'h5687] = 8'h4C;
mem[16'h5688] = 8'h03;
mem[16'h5689] = 8'h40;
mem[16'h568A] = 8'h00;
mem[16'h568B] = 8'h52;
mem[16'h568C] = 8'h03;
mem[16'h568D] = 8'h40;
mem[16'h568E] = 8'h00;
mem[16'h568F] = 8'h12;
mem[16'h5690] = 8'h04;
mem[16'h5691] = 8'h40;
mem[16'h5692] = 8'h00;
mem[16'h5693] = 8'h12;
mem[16'h5694] = 8'h04;
mem[16'h5695] = 8'h40;
mem[16'h5696] = 8'h00;
mem[16'h5697] = 8'h52;
mem[16'h5698] = 8'h03;
mem[16'h5699] = 8'h40;
mem[16'h569A] = 8'h00;
mem[16'h569B] = 8'h4C;
mem[16'h569C] = 8'h03;
mem[16'h569D] = 8'h40;
mem[16'h569E] = 8'h00;
mem[16'h569F] = 8'h00;
mem[16'h56A0] = 8'h1E;
mem[16'h56A1] = 8'h78;
mem[16'h56A2] = 8'h00;
mem[16'h56A3] = 8'h00;
mem[16'h56A4] = 8'h3C;
mem[16'h56A5] = 8'h70;
mem[16'h56A6] = 8'h01;
mem[16'h56A7] = 8'h18;
mem[16'h56A8] = 8'h07;
mem[16'h56A9] = 8'h00;
mem[16'h56AA] = 8'h01;
mem[16'h56AB] = 8'h24;
mem[16'h56AC] = 8'h07;
mem[16'h56AD] = 8'h00;
mem[16'h56AE] = 8'h01;
mem[16'h56AF] = 8'h24;
mem[16'h56B0] = 8'h08;
mem[16'h56B1] = 8'h00;
mem[16'h56B2] = 8'h01;
mem[16'h56B3] = 8'h24;
mem[16'h56B4] = 8'h08;
mem[16'h56B5] = 8'h00;
mem[16'h56B6] = 8'h01;
mem[16'h56B7] = 8'h24;
mem[16'h56B8] = 8'h07;
mem[16'h56B9] = 8'h00;
mem[16'h56BA] = 8'h01;
mem[16'h56BB] = 8'h18;
mem[16'h56BC] = 8'h07;
mem[16'h56BD] = 8'h00;
mem[16'h56BE] = 8'h01;
mem[16'h56BF] = 8'h00;
mem[16'h56C0] = 8'h3C;
mem[16'h56C1] = 8'h70;
mem[16'h56C2] = 8'h01;
mem[16'h56C3] = 8'h00;
mem[16'h56C4] = 8'h78;
mem[16'h56C5] = 8'h60;
mem[16'h56C6] = 8'h03;
mem[16'h56C7] = 8'h30;
mem[16'h56C8] = 8'h0E;
mem[16'h56C9] = 8'h00;
mem[16'h56CA] = 8'h02;
mem[16'h56CB] = 8'h48;
mem[16'h56CC] = 8'h0E;
mem[16'h56CD] = 8'h00;
mem[16'h56CE] = 8'h02;
mem[16'h56CF] = 8'h48;
mem[16'h56D0] = 8'h10;
mem[16'h56D1] = 8'h00;
mem[16'h56D2] = 8'h02;
mem[16'h56D3] = 8'h48;
mem[16'h56D4] = 8'h10;
mem[16'h56D5] = 8'h00;
mem[16'h56D6] = 8'h02;
mem[16'h56D7] = 8'h48;
mem[16'h56D8] = 8'h0E;
mem[16'h56D9] = 8'h00;
mem[16'h56DA] = 8'h02;
mem[16'h56DB] = 8'h30;
mem[16'h56DC] = 8'h0E;
mem[16'h56DD] = 8'h00;
mem[16'h56DE] = 8'h02;
mem[16'h56DF] = 8'h00;
mem[16'h56E0] = 8'h78;
mem[16'h56E1] = 8'h60;
mem[16'h56E2] = 8'h03;
mem[16'h56E3] = 8'h00;
mem[16'h56E4] = 8'h70;
mem[16'h56E5] = 8'h41;
mem[16'h56E6] = 8'h07;
mem[16'h56E7] = 8'h60;
mem[16'h56E8] = 8'h1C;
mem[16'h56E9] = 8'h00;
mem[16'h56EA] = 8'h04;
mem[16'h56EB] = 8'h10;
mem[16'h56EC] = 8'h1D;
mem[16'h56ED] = 8'h00;
mem[16'h56EE] = 8'h04;
mem[16'h56EF] = 8'h10;
mem[16'h56F0] = 8'h21;
mem[16'h56F1] = 8'h00;
mem[16'h56F2] = 8'h04;
mem[16'h56F3] = 8'h10;
mem[16'h56F4] = 8'h21;
mem[16'h56F5] = 8'h00;
mem[16'h56F6] = 8'h04;
mem[16'h56F7] = 8'h10;
mem[16'h56F8] = 8'h1D;
mem[16'h56F9] = 8'h00;
mem[16'h56FA] = 8'h04;
mem[16'h56FB] = 8'h60;
mem[16'h56FC] = 8'h1C;
mem[16'h56FD] = 8'h00;
mem[16'h56FE] = 8'h04;
mem[16'h56FF] = 8'h00;
mem[16'h5700] = 8'h70;
mem[16'h5701] = 8'h41;
mem[16'h5702] = 8'h07;
mem[16'h5703] = 8'h00;
mem[16'h5704] = 8'h60;
mem[16'h5705] = 8'h03;
mem[16'h5706] = 8'h0F;
mem[16'h5707] = 8'h40;
mem[16'h5708] = 8'h39;
mem[16'h5709] = 8'h00;
mem[16'h570A] = 8'h08;
mem[16'h570B] = 8'h20;
mem[16'h570C] = 8'h3A;
mem[16'h570D] = 8'h00;
mem[16'h570E] = 8'h08;
mem[16'h570F] = 8'h20;
mem[16'h5710] = 8'h42;
mem[16'h5711] = 8'h00;
mem[16'h5712] = 8'h08;
mem[16'h5713] = 8'h20;
mem[16'h5714] = 8'h42;
mem[16'h5715] = 8'h00;
mem[16'h5716] = 8'h08;
mem[16'h5717] = 8'h20;
mem[16'h5718] = 8'h3A;
mem[16'h5719] = 8'h00;
mem[16'h571A] = 8'h08;
mem[16'h571B] = 8'h40;
mem[16'h571C] = 8'h39;
mem[16'h571D] = 8'h00;
mem[16'h571E] = 8'h08;
mem[16'h571F] = 8'h00;
mem[16'h5720] = 8'h60;
mem[16'h5721] = 8'h03;
mem[16'h5722] = 8'h0F;
mem[16'h5723] = 8'h00;
mem[16'h5724] = 8'h40;
mem[16'h5725] = 8'h07;
mem[16'h5726] = 8'h1E;
mem[16'h5727] = 8'h00;
mem[16'h5728] = 8'h73;
mem[16'h5729] = 8'h00;
mem[16'h572A] = 8'h10;
mem[16'h572B] = 8'h40;
mem[16'h572C] = 8'h74;
mem[16'h572D] = 8'h00;
mem[16'h572E] = 8'h10;
mem[16'h572F] = 8'h40;
mem[16'h5730] = 8'h04;
mem[16'h5731] = 8'h01;
mem[16'h5732] = 8'h10;
mem[16'h5733] = 8'h40;
mem[16'h5734] = 8'h04;
mem[16'h5735] = 8'h01;
mem[16'h5736] = 8'h10;
mem[16'h5737] = 8'h40;
mem[16'h5738] = 8'h74;
mem[16'h5739] = 8'h00;
mem[16'h573A] = 8'h10;
mem[16'h573B] = 8'h00;
mem[16'h573C] = 8'h73;
mem[16'h573D] = 8'h00;
mem[16'h573E] = 8'h10;
mem[16'h573F] = 8'h00;
mem[16'h5740] = 8'h40;
mem[16'h5741] = 8'h07;
mem[16'h5742] = 8'h1E;
mem[16'h5743] = 8'hAE;
mem[16'h5744] = 8'hAB;
mem[16'h5745] = 8'h4A;
mem[16'h5746] = 8'hCA;
mem[16'h5747] = 8'h30;
mem[16'h5748] = 8'h29;
mem[16'h5749] = 8'h86;
mem[16'h574A] = 8'h70;
mem[16'h574B] = 8'hBD;
mem[16'h574C] = 8'hEB;
mem[16'h574D] = 8'h60;
mem[16'h574E] = 8'hC9;
mem[16'h574F] = 8'h02;
mem[16'h5750] = 8'h90;
mem[16'h5751] = 8'h0E;
mem[16'h5752] = 8'h38;
mem[16'h5753] = 8'hE9;
mem[16'h5754] = 8'h02;
mem[16'h5755] = 8'h9D;
mem[16'h5756] = 8'hEB;
mem[16'h5757] = 8'h60;
mem[16'h5758] = 8'h20;
mem[16'h5759] = 8'h73;
mem[16'h575A] = 8'h57;
mem[16'h575B] = 8'hA6;
mem[16'h575C] = 8'h70;
mem[16'h575D] = 8'h4C;
mem[16'h575E] = 8'h46;
mem[16'h575F] = 8'h57;
mem[16'h5760] = 8'h20;
mem[16'h5761] = 8'hB7;
mem[16'h5762] = 8'h60;
mem[16'h5763] = 8'hA6;
mem[16'h5764] = 8'h70;
mem[16'h5765] = 8'hA9;
mem[16'h5766] = 8'hFE;
mem[16'h5767] = 8'h9D;
mem[16'h5768] = 8'hEB;
mem[16'h5769] = 8'h60;
mem[16'h576A] = 8'h20;
mem[16'h576B] = 8'hB7;
mem[16'h576C] = 8'h60;
mem[16'h576D] = 8'hA6;
mem[16'h576E] = 8'h70;
mem[16'h576F] = 8'h4C;
mem[16'h5770] = 8'h46;
mem[16'h5771] = 8'h57;
mem[16'h5772] = 8'h60;
mem[16'h5773] = 8'hA6;
mem[16'h5774] = 8'h70;
mem[16'h5775] = 8'hBD;
mem[16'h5776] = 8'hEF;
mem[16'h5777] = 8'h60;
mem[16'h5778] = 8'h85;
mem[16'h5779] = 8'h56;
mem[16'h577A] = 8'hBC;
mem[16'h577B] = 8'hEB;
mem[16'h577C] = 8'h60;
mem[16'h577D] = 8'h84;
mem[16'h577E] = 8'h57;
mem[16'h577F] = 8'hB9;
mem[16'h5780] = 8'h3E;
mem[16'h5781] = 8'h8C;
mem[16'h5782] = 8'hAA;
mem[16'h5783] = 8'hBD;
mem[16'h5784] = 8'h94;
mem[16'h5785] = 8'h8E;
mem[16'h5786] = 8'hAA;
mem[16'h5787] = 8'hBD;
mem[16'h5788] = 8'h99;
mem[16'h5789] = 8'h57;
mem[16'h578A] = 8'hBC;
mem[16'h578B] = 8'hA0;
mem[16'h578C] = 8'h57;
mem[16'h578D] = 8'h20;
mem[16'h578E] = 8'hD1;
mem[16'h578F] = 8'h8A;
mem[16'h5790] = 8'hA9;
mem[16'h5791] = 8'h20;
mem[16'h5792] = 8'h8D;
mem[16'h5793] = 8'hCA;
mem[16'h5794] = 8'h8A;
mem[16'h5795] = 8'h20;
mem[16'h5796] = 8'h79;
mem[16'h5797] = 8'h8A;
mem[16'h5798] = 8'h60;
mem[16'h5799] = 8'hA7;
mem[16'h579A] = 8'hC7;
mem[16'h579B] = 8'hE7;
mem[16'h579C] = 8'h07;
mem[16'h579D] = 8'h27;
mem[16'h579E] = 8'h47;
mem[16'h579F] = 8'h67;
mem[16'h57A0] = 8'h57;
mem[16'h57A1] = 8'h57;
mem[16'h57A2] = 8'h57;
mem[16'h57A3] = 8'h58;
mem[16'h57A4] = 8'h58;
mem[16'h57A5] = 8'h58;
mem[16'h57A6] = 8'h58;
mem[16'h57A7] = 8'h18;
mem[16'h57A8] = 8'h73;
mem[16'h57A9] = 8'h04;
mem[16'h57AA] = 8'h00;
mem[16'h57AB] = 8'h04;
mem[16'h57AC] = 8'h00;
mem[16'h57AD] = 8'h0E;
mem[16'h57AE] = 8'h00;
mem[16'h57AF] = 8'h0E;
mem[16'h57B0] = 8'h00;
mem[16'h57B1] = 8'h32;
mem[16'h57B2] = 8'h00;
mem[16'h57B3] = 8'h01;
mem[16'h57B4] = 8'h0A;
mem[16'h57B5] = 8'h0E;
mem[16'h57B6] = 8'h00;
mem[16'h57B7] = 8'h01;
mem[16'h57B8] = 8'h0A;
mem[16'h57B9] = 8'h0E;
mem[16'h57BA] = 8'h00;
mem[16'h57BB] = 8'h0E;
mem[16'h57BC] = 8'h00;
mem[16'h57BD] = 8'h32;
mem[16'h57BE] = 8'h00;
mem[16'h57BF] = 8'h04;
mem[16'h57C0] = 8'h00;
mem[16'h57C1] = 8'h0E;
mem[16'h57C2] = 8'h00;
mem[16'h57C3] = 8'h18;
mem[16'h57C4] = 8'h73;
mem[16'h57C5] = 8'h04;
mem[16'h57C6] = 8'h00;
mem[16'h57C7] = 8'h30;
mem[16'h57C8] = 8'h66;
mem[16'h57C9] = 8'h09;
mem[16'h57CA] = 8'h00;
mem[16'h57CB] = 8'h08;
mem[16'h57CC] = 8'h00;
mem[16'h57CD] = 8'h1C;
mem[16'h57CE] = 8'h00;
mem[16'h57CF] = 8'h1C;
mem[16'h57D0] = 8'h00;
mem[16'h57D1] = 8'h64;
mem[16'h57D2] = 8'h00;
mem[16'h57D3] = 8'h02;
mem[16'h57D4] = 8'h14;
mem[16'h57D5] = 8'h1C;
mem[16'h57D6] = 8'h00;
mem[16'h57D7] = 8'h02;
mem[16'h57D8] = 8'h14;
mem[16'h57D9] = 8'h1C;
mem[16'h57DA] = 8'h00;
mem[16'h57DB] = 8'h1C;
mem[16'h57DC] = 8'h00;
mem[16'h57DD] = 8'h64;
mem[16'h57DE] = 8'h00;
mem[16'h57DF] = 8'h08;
mem[16'h57E0] = 8'h00;
mem[16'h57E1] = 8'h1C;
mem[16'h57E2] = 8'h00;
mem[16'h57E3] = 8'h30;
mem[16'h57E4] = 8'h66;
mem[16'h57E5] = 8'h09;
mem[16'h57E6] = 8'h00;
mem[16'h57E7] = 8'h60;
mem[16'h57E8] = 8'h4C;
mem[16'h57E9] = 8'h13;
mem[16'h57EA] = 8'h00;
mem[16'h57EB] = 8'h10;
mem[16'h57EC] = 8'h00;
mem[16'h57ED] = 8'h38;
mem[16'h57EE] = 8'h00;
mem[16'h57EF] = 8'h38;
mem[16'h57F0] = 8'h00;
mem[16'h57F1] = 8'h48;
mem[16'h57F2] = 8'h01;
mem[16'h57F3] = 8'h04;
mem[16'h57F4] = 8'h28;
mem[16'h57F5] = 8'h38;
mem[16'h57F6] = 8'h00;
mem[16'h57F7] = 8'h04;
mem[16'h57F8] = 8'h28;
mem[16'h57F9] = 8'h38;
mem[16'h57FA] = 8'h00;
mem[16'h57FB] = 8'h38;
mem[16'h57FC] = 8'h00;
mem[16'h57FD] = 8'h48;
mem[16'h57FE] = 8'h01;
mem[16'h57FF] = 8'h10;
mem[16'h5800] = 8'h00;
mem[16'h5801] = 8'h38;
mem[16'h5802] = 8'h00;
mem[16'h5803] = 8'h60;
mem[16'h5804] = 8'h4C;
mem[16'h5805] = 8'h13;
mem[16'h5806] = 8'h00;
mem[16'h5807] = 8'h40;
mem[16'h5808] = 8'h19;
mem[16'h5809] = 8'h27;
mem[16'h580A] = 8'h00;
mem[16'h580B] = 8'h20;
mem[16'h580C] = 8'h00;
mem[16'h580D] = 8'h70;
mem[16'h580E] = 8'h00;
mem[16'h580F] = 8'h70;
mem[16'h5810] = 8'h00;
mem[16'h5811] = 8'h10;
mem[16'h5812] = 8'h03;
mem[16'h5813] = 8'h08;
mem[16'h5814] = 8'h50;
mem[16'h5815] = 8'h70;
mem[16'h5816] = 8'h00;
mem[16'h5817] = 8'h08;
mem[16'h5818] = 8'h50;
mem[16'h5819] = 8'h70;
mem[16'h581A] = 8'h00;
mem[16'h581B] = 8'h70;
mem[16'h581C] = 8'h00;
mem[16'h581D] = 8'h10;
mem[16'h581E] = 8'h03;
mem[16'h581F] = 8'h20;
mem[16'h5820] = 8'h00;
mem[16'h5821] = 8'h70;
mem[16'h5822] = 8'h00;
mem[16'h5823] = 8'h40;
mem[16'h5824] = 8'h19;
mem[16'h5825] = 8'h27;
mem[16'h5826] = 8'h00;
mem[16'h5827] = 8'h00;
mem[16'h5828] = 8'h33;
mem[16'h5829] = 8'h4E;
mem[16'h582A] = 8'h00;
mem[16'h582B] = 8'h40;
mem[16'h582C] = 8'h00;
mem[16'h582D] = 8'h60;
mem[16'h582E] = 8'h01;
mem[16'h582F] = 8'h60;
mem[16'h5830] = 8'h01;
mem[16'h5831] = 8'h20;
mem[16'h5832] = 8'h06;
mem[16'h5833] = 8'h10;
mem[16'h5834] = 8'h20;
mem[16'h5835] = 8'h61;
mem[16'h5836] = 8'h01;
mem[16'h5837] = 8'h10;
mem[16'h5838] = 8'h20;
mem[16'h5839] = 8'h61;
mem[16'h583A] = 8'h01;
mem[16'h583B] = 8'h60;
mem[16'h583C] = 8'h01;
mem[16'h583D] = 8'h20;
mem[16'h583E] = 8'h06;
mem[16'h583F] = 8'h40;
mem[16'h5840] = 8'h00;
mem[16'h5841] = 8'h60;
mem[16'h5842] = 8'h01;
mem[16'h5843] = 8'h00;
mem[16'h5844] = 8'h33;
mem[16'h5845] = 8'h4E;
mem[16'h5846] = 8'h00;
mem[16'h5847] = 8'h00;
mem[16'h5848] = 8'h66;
mem[16'h5849] = 8'h1C;
mem[16'h584A] = 8'h01;
mem[16'h584B] = 8'h00;
mem[16'h584C] = 8'h01;
mem[16'h584D] = 8'h40;
mem[16'h584E] = 8'h03;
mem[16'h584F] = 8'h40;
mem[16'h5850] = 8'h03;
mem[16'h5851] = 8'h40;
mem[16'h5852] = 8'h0C;
mem[16'h5853] = 8'h20;
mem[16'h5854] = 8'h40;
mem[16'h5855] = 8'h42;
mem[16'h5856] = 8'h03;
mem[16'h5857] = 8'h20;
mem[16'h5858] = 8'h40;
mem[16'h5859] = 8'h42;
mem[16'h585A] = 8'h03;
mem[16'h585B] = 8'h40;
mem[16'h585C] = 8'h03;
mem[16'h585D] = 8'h40;
mem[16'h585E] = 8'h0C;
mem[16'h585F] = 8'h00;
mem[16'h5860] = 8'h01;
mem[16'h5861] = 8'h40;
mem[16'h5862] = 8'h03;
mem[16'h5863] = 8'h00;
mem[16'h5864] = 8'h66;
mem[16'h5865] = 8'h1C;
mem[16'h5866] = 8'h01;
mem[16'h5867] = 8'h00;
mem[16'h5868] = 8'h4C;
mem[16'h5869] = 8'h39;
mem[16'h586A] = 8'h02;
mem[16'h586B] = 8'h00;
mem[16'h586C] = 8'h02;
mem[16'h586D] = 8'h00;
mem[16'h586E] = 8'h07;
mem[16'h586F] = 8'h00;
mem[16'h5870] = 8'h07;
mem[16'h5871] = 8'h00;
mem[16'h5872] = 8'h19;
mem[16'h5873] = 8'h40;
mem[16'h5874] = 8'h00;
mem[16'h5875] = 8'h05;
mem[16'h5876] = 8'h07;
mem[16'h5877] = 8'h40;
mem[16'h5878] = 8'h00;
mem[16'h5879] = 8'h05;
mem[16'h587A] = 8'h07;
mem[16'h587B] = 8'h00;
mem[16'h587C] = 8'h07;
mem[16'h587D] = 8'h00;
mem[16'h587E] = 8'h19;
mem[16'h587F] = 8'h00;
mem[16'h5880] = 8'h02;
mem[16'h5881] = 8'h00;
mem[16'h5882] = 8'h07;
mem[16'h5883] = 8'h00;
mem[16'h5884] = 8'h4C;
mem[16'h5885] = 8'h39;
mem[16'h5886] = 8'h02;
mem[16'h5887] = 8'hAE;
mem[16'h5888] = 8'hAC;
mem[16'h5889] = 8'h4A;
mem[16'h588A] = 8'hCA;
mem[16'h588B] = 8'h30;
mem[16'h588C] = 8'h29;
mem[16'h588D] = 8'h86;
mem[16'h588E] = 8'h70;
mem[16'h588F] = 8'hBD;
mem[16'h5890] = 8'h2A;
mem[16'h5891] = 8'h61;
mem[16'h5892] = 8'hC9;
mem[16'h5893] = 8'h02;
mem[16'h5894] = 8'h90;
mem[16'h5895] = 8'h0E;
mem[16'h5896] = 8'h38;
mem[16'h5897] = 8'hE9;
mem[16'h5898] = 8'h02;
mem[16'h5899] = 8'h9D;
mem[16'h589A] = 8'h2A;
mem[16'h589B] = 8'h61;
mem[16'h589C] = 8'h20;
mem[16'h589D] = 8'hB7;
mem[16'h589E] = 8'h58;
mem[16'h589F] = 8'hA6;
mem[16'h58A0] = 8'h70;
mem[16'h58A1] = 8'h4C;
mem[16'h58A2] = 8'h8A;
mem[16'h58A3] = 8'h58;
mem[16'h58A4] = 8'h20;
mem[16'h58A5] = 8'hF3;
mem[16'h58A6] = 8'h60;
mem[16'h58A7] = 8'hA6;
mem[16'h58A8] = 8'h70;
mem[16'h58A9] = 8'hA9;
mem[16'h58AA] = 8'hFE;
mem[16'h58AB] = 8'h9D;
mem[16'h58AC] = 8'h2A;
mem[16'h58AD] = 8'h61;
mem[16'h58AE] = 8'h20;
mem[16'h58AF] = 8'hF3;
mem[16'h58B0] = 8'h60;
mem[16'h58B1] = 8'hA6;
mem[16'h58B2] = 8'h70;
mem[16'h58B3] = 8'h4C;
mem[16'h58B4] = 8'h8A;
mem[16'h58B5] = 8'h58;
mem[16'h58B6] = 8'h60;
mem[16'h58B7] = 8'hA6;
mem[16'h58B8] = 8'h70;
mem[16'h58B9] = 8'hBD;
mem[16'h58BA] = 8'h2E;
mem[16'h58BB] = 8'h61;
mem[16'h58BC] = 8'h85;
mem[16'h58BD] = 8'h56;
mem[16'h58BE] = 8'hBC;
mem[16'h58BF] = 8'h2A;
mem[16'h58C0] = 8'h61;
mem[16'h58C1] = 8'h84;
mem[16'h58C2] = 8'h57;
mem[16'h58C3] = 8'hB9;
mem[16'h58C4] = 8'h3E;
mem[16'h58C5] = 8'h8C;
mem[16'h58C6] = 8'hAA;
mem[16'h58C7] = 8'hBD;
mem[16'h58C8] = 8'h94;
mem[16'h58C9] = 8'h8E;
mem[16'h58CA] = 8'hAA;
mem[16'h58CB] = 8'hBD;
mem[16'h58CC] = 8'hDD;
mem[16'h58CD] = 8'h58;
mem[16'h58CE] = 8'hBC;
mem[16'h58CF] = 8'hE4;
mem[16'h58D0] = 8'h58;
mem[16'h58D1] = 8'h20;
mem[16'h58D2] = 8'hD1;
mem[16'h58D3] = 8'h8A;
mem[16'h58D4] = 8'hA9;
mem[16'h58D5] = 8'h24;
mem[16'h58D6] = 8'h8D;
mem[16'h58D7] = 8'hCA;
mem[16'h58D8] = 8'h8A;
mem[16'h58D9] = 8'h20;
mem[16'h58DA] = 8'h79;
mem[16'h58DB] = 8'h8A;
mem[16'h58DC] = 8'h60;
mem[16'h58DD] = 8'hEB;
mem[16'h58DE] = 8'h0F;
mem[16'h58DF] = 8'h33;
mem[16'h58E0] = 8'h57;
mem[16'h58E1] = 8'h7B;
mem[16'h58E2] = 8'h9F;
mem[16'h58E3] = 8'hC3;
mem[16'h58E4] = 8'h58;
mem[16'h58E5] = 8'h59;
mem[16'h58E6] = 8'h59;
mem[16'h58E7] = 8'h59;
mem[16'h58E8] = 8'h59;
mem[16'h58E9] = 8'h59;
mem[16'h58EA] = 8'h59;
mem[16'h58EB] = 8'h33;
mem[16'h58EC] = 8'h40;
mem[16'h58ED] = 8'h19;
mem[16'h58EE] = 8'h00;
mem[16'h58EF] = 8'h73;
mem[16'h58F0] = 8'h60;
mem[16'h58F1] = 8'h19;
mem[16'h58F2] = 8'h00;
mem[16'h58F3] = 8'h0E;
mem[16'h58F4] = 8'h00;
mem[16'h58F5] = 8'h0E;
mem[16'h58F6] = 8'h00;
mem[16'h58F7] = 8'h41;
mem[16'h58F8] = 8'h08;
mem[16'h58F9] = 8'h68;
mem[16'h58FA] = 8'h00;
mem[16'h58FB] = 8'h41;
mem[16'h58FC] = 8'h08;
mem[16'h58FD] = 8'h04;
mem[16'h58FE] = 8'h00;
mem[16'h58FF] = 8'h41;
mem[16'h5900] = 8'h08;
mem[16'h5901] = 8'h68;
mem[16'h5902] = 8'h00;
mem[16'h5903] = 8'h0E;
mem[16'h5904] = 8'h00;
mem[16'h5905] = 8'h0E;
mem[16'h5906] = 8'h00;
mem[16'h5907] = 8'h73;
mem[16'h5908] = 8'h60;
mem[16'h5909] = 8'h19;
mem[16'h590A] = 8'h00;
mem[16'h590B] = 8'h33;
mem[16'h590C] = 8'h40;
mem[16'h590D] = 8'h19;
mem[16'h590E] = 8'h00;
mem[16'h590F] = 8'h66;
mem[16'h5910] = 8'h00;
mem[16'h5911] = 8'h33;
mem[16'h5912] = 8'h00;
mem[16'h5913] = 8'h66;
mem[16'h5914] = 8'h41;
mem[16'h5915] = 8'h33;
mem[16'h5916] = 8'h00;
mem[16'h5917] = 8'h1C;
mem[16'h5918] = 8'h00;
mem[16'h5919] = 8'h1C;
mem[16'h591A] = 8'h00;
mem[16'h591B] = 8'h02;
mem[16'h591C] = 8'h11;
mem[16'h591D] = 8'h50;
mem[16'h591E] = 8'h01;
mem[16'h591F] = 8'h02;
mem[16'h5920] = 8'h11;
mem[16'h5921] = 8'h08;
mem[16'h5922] = 8'h00;
mem[16'h5923] = 8'h02;
mem[16'h5924] = 8'h11;
mem[16'h5925] = 8'h50;
mem[16'h5926] = 8'h01;
mem[16'h5927] = 8'h1C;
mem[16'h5928] = 8'h00;
mem[16'h5929] = 8'h1C;
mem[16'h592A] = 8'h00;
mem[16'h592B] = 8'h66;
mem[16'h592C] = 8'h41;
mem[16'h592D] = 8'h33;
mem[16'h592E] = 8'h00;
mem[16'h592F] = 8'h66;
mem[16'h5930] = 8'h00;
mem[16'h5931] = 8'h33;
mem[16'h5932] = 8'h00;
mem[16'h5933] = 8'h4C;
mem[16'h5934] = 8'h01;
mem[16'h5935] = 8'h66;
mem[16'h5936] = 8'h00;
mem[16'h5937] = 8'h4C;
mem[16'h5938] = 8'h03;
mem[16'h5939] = 8'h67;
mem[16'h593A] = 8'h00;
mem[16'h593B] = 8'h38;
mem[16'h593C] = 8'h00;
mem[16'h593D] = 8'h38;
mem[16'h593E] = 8'h00;
mem[16'h593F] = 8'h04;
mem[16'h5940] = 8'h22;
mem[16'h5941] = 8'h20;
mem[16'h5942] = 8'h03;
mem[16'h5943] = 8'h04;
mem[16'h5944] = 8'h22;
mem[16'h5945] = 8'h10;
mem[16'h5946] = 8'h00;
mem[16'h5947] = 8'h04;
mem[16'h5948] = 8'h22;
mem[16'h5949] = 8'h20;
mem[16'h594A] = 8'h03;
mem[16'h594B] = 8'h38;
mem[16'h594C] = 8'h00;
mem[16'h594D] = 8'h38;
mem[16'h594E] = 8'h00;
mem[16'h594F] = 8'h4C;
mem[16'h5950] = 8'h03;
mem[16'h5951] = 8'h67;
mem[16'h5952] = 8'h00;
mem[16'h5953] = 8'h4C;
mem[16'h5954] = 8'h01;
mem[16'h5955] = 8'h66;
mem[16'h5956] = 8'h00;
mem[16'h5957] = 8'h18;
mem[16'h5958] = 8'h03;
mem[16'h5959] = 8'h4C;
mem[16'h595A] = 8'h01;
mem[16'h595B] = 8'h18;
mem[16'h595C] = 8'h07;
mem[16'h595D] = 8'h4E;
mem[16'h595E] = 8'h01;
mem[16'h595F] = 8'h70;
mem[16'h5960] = 8'h00;
mem[16'h5961] = 8'h70;
mem[16'h5962] = 8'h00;
mem[16'h5963] = 8'h08;
mem[16'h5964] = 8'h44;
mem[16'h5965] = 8'h40;
mem[16'h5966] = 8'h06;
mem[16'h5967] = 8'h08;
mem[16'h5968] = 8'h44;
mem[16'h5969] = 8'h20;
mem[16'h596A] = 8'h00;
mem[16'h596B] = 8'h08;
mem[16'h596C] = 8'h44;
mem[16'h596D] = 8'h40;
mem[16'h596E] = 8'h06;
mem[16'h596F] = 8'h70;
mem[16'h5970] = 8'h00;
mem[16'h5971] = 8'h70;
mem[16'h5972] = 8'h00;
mem[16'h5973] = 8'h18;
mem[16'h5974] = 8'h07;
mem[16'h5975] = 8'h4E;
mem[16'h5976] = 8'h01;
mem[16'h5977] = 8'h18;
mem[16'h5978] = 8'h03;
mem[16'h5979] = 8'h4C;
mem[16'h597A] = 8'h01;
mem[16'h597B] = 8'h30;
mem[16'h597C] = 8'h06;
mem[16'h597D] = 8'h18;
mem[16'h597E] = 8'h03;
mem[16'h597F] = 8'h30;
mem[16'h5980] = 8'h0E;
mem[16'h5981] = 8'h1C;
mem[16'h5982] = 8'h03;
mem[16'h5983] = 8'h60;
mem[16'h5984] = 8'h01;
mem[16'h5985] = 8'h60;
mem[16'h5986] = 8'h01;
mem[16'h5987] = 8'h10;
mem[16'h5988] = 8'h08;
mem[16'h5989] = 8'h01;
mem[16'h598A] = 8'h0D;
mem[16'h598B] = 8'h10;
mem[16'h598C] = 8'h08;
mem[16'h598D] = 8'h41;
mem[16'h598E] = 8'h00;
mem[16'h598F] = 8'h10;
mem[16'h5990] = 8'h08;
mem[16'h5991] = 8'h01;
mem[16'h5992] = 8'h0D;
mem[16'h5993] = 8'h60;
mem[16'h5994] = 8'h01;
mem[16'h5995] = 8'h60;
mem[16'h5996] = 8'h01;
mem[16'h5997] = 8'h30;
mem[16'h5998] = 8'h0E;
mem[16'h5999] = 8'h1C;
mem[16'h599A] = 8'h03;
mem[16'h599B] = 8'h30;
mem[16'h599C] = 8'h06;
mem[16'h599D] = 8'h18;
mem[16'h599E] = 8'h03;
mem[16'h599F] = 8'h60;
mem[16'h59A0] = 8'h0C;
mem[16'h59A1] = 8'h30;
mem[16'h59A2] = 8'h06;
mem[16'h59A3] = 8'h60;
mem[16'h59A4] = 8'h1C;
mem[16'h59A5] = 8'h38;
mem[16'h59A6] = 8'h06;
mem[16'h59A7] = 8'h40;
mem[16'h59A8] = 8'h03;
mem[16'h59A9] = 8'h40;
mem[16'h59AA] = 8'h03;
mem[16'h59AB] = 8'h20;
mem[16'h59AC] = 8'h10;
mem[16'h59AD] = 8'h02;
mem[16'h59AE] = 8'h1A;
mem[16'h59AF] = 8'h20;
mem[16'h59B0] = 8'h10;
mem[16'h59B1] = 8'h02;
mem[16'h59B2] = 8'h01;
mem[16'h59B3] = 8'h20;
mem[16'h59B4] = 8'h10;
mem[16'h59B5] = 8'h02;
mem[16'h59B6] = 8'h1A;
mem[16'h59B7] = 8'h40;
mem[16'h59B8] = 8'h03;
mem[16'h59B9] = 8'h40;
mem[16'h59BA] = 8'h03;
mem[16'h59BB] = 8'h60;
mem[16'h59BC] = 8'h1C;
mem[16'h59BD] = 8'h38;
mem[16'h59BE] = 8'h06;
mem[16'h59BF] = 8'h60;
mem[16'h59C0] = 8'h0C;
mem[16'h59C1] = 8'h30;
mem[16'h59C2] = 8'h06;
mem[16'h59C3] = 8'h40;
mem[16'h59C4] = 8'h19;
mem[16'h59C5] = 8'h60;
mem[16'h59C6] = 8'h0C;
mem[16'h59C7] = 8'h40;
mem[16'h59C8] = 8'h39;
mem[16'h59C9] = 8'h70;
mem[16'h59CA] = 8'h0C;
mem[16'h59CB] = 8'h00;
mem[16'h59CC] = 8'h07;
mem[16'h59CD] = 8'h00;
mem[16'h59CE] = 8'h07;
mem[16'h59CF] = 8'h40;
mem[16'h59D0] = 8'h20;
mem[16'h59D1] = 8'h04;
mem[16'h59D2] = 8'h34;
mem[16'h59D3] = 8'h40;
mem[16'h59D4] = 8'h20;
mem[16'h59D5] = 8'h04;
mem[16'h59D6] = 8'h02;
mem[16'h59D7] = 8'h40;
mem[16'h59D8] = 8'h20;
mem[16'h59D9] = 8'h04;
mem[16'h59DA] = 8'h34;
mem[16'h59DB] = 8'h00;
mem[16'h59DC] = 8'h07;
mem[16'h59DD] = 8'h00;
mem[16'h59DE] = 8'h07;
mem[16'h59DF] = 8'h40;
mem[16'h59E0] = 8'h39;
mem[16'h59E1] = 8'h70;
mem[16'h59E2] = 8'h0C;
mem[16'h59E3] = 8'h40;
mem[16'h59E4] = 8'h19;
mem[16'h59E5] = 8'h60;
mem[16'h59E6] = 8'h0C;
mem[16'h59E7] = 8'hAE;
mem[16'h59E8] = 8'hB0;
mem[16'h59E9] = 8'h4A;
mem[16'h59EA] = 8'hCA;
mem[16'h59EB] = 8'hE0;
mem[16'h59EC] = 8'h08;
mem[16'h59ED] = 8'h90;
mem[16'h59EE] = 8'h2E;
mem[16'h59EF] = 8'h86;
mem[16'h59F0] = 8'h70;
mem[16'h59F1] = 8'hBD;
mem[16'h59F2] = 8'h75;
mem[16'h59F3] = 8'h5B;
mem[16'h59F4] = 8'hD0;
mem[16'h59F5] = 8'h28;
mem[16'h59F6] = 8'hBD;
mem[16'h59F7] = 8'h2C;
mem[16'h59F8] = 8'h5F;
mem[16'h59F9] = 8'hC9;
mem[16'h59FA] = 8'h02;
mem[16'h59FB] = 8'h90;
mem[16'h59FC] = 8'h0E;
mem[16'h59FD] = 8'h38;
mem[16'h59FE] = 8'hE9;
mem[16'h59FF] = 8'h02;
mem[16'h5A00] = 8'h9D;
mem[16'h5A01] = 8'h2C;
mem[16'h5A02] = 8'h5F;
mem[16'h5A03] = 8'h20;
mem[16'h5A04] = 8'h91;
mem[16'h5A05] = 8'h5B;
mem[16'h5A06] = 8'hA6;
mem[16'h5A07] = 8'h70;
mem[16'h5A08] = 8'h4C;
mem[16'h5A09] = 8'hEA;
mem[16'h5A0A] = 8'h59;
mem[16'h5A0B] = 8'h20;
mem[16'h5A0C] = 8'hC4;
mem[16'h5A0D] = 8'h72;
mem[16'h5A0E] = 8'hA6;
mem[16'h5A0F] = 8'h70;
mem[16'h5A10] = 8'hA9;
mem[16'h5A11] = 8'hEB;
mem[16'h5A12] = 8'h9D;
mem[16'h5A13] = 8'h2C;
mem[16'h5A14] = 8'h5F;
mem[16'h5A15] = 8'h20;
mem[16'h5A16] = 8'hC4;
mem[16'h5A17] = 8'h72;
mem[16'h5A18] = 8'hA6;
mem[16'h5A19] = 8'h70;
mem[16'h5A1A] = 8'h4C;
mem[16'h5A1B] = 8'hEA;
mem[16'h5A1C] = 8'h59;
mem[16'h5A1D] = 8'h60;
mem[16'h5A1E] = 8'hC9;
mem[16'h5A1F] = 8'h24;
mem[16'h5A20] = 8'hD0;
mem[16'h5A21] = 8'h05;
mem[16'h5A22] = 8'h20;
mem[16'h5A23] = 8'hB1;
mem[16'h5A24] = 8'h75;
mem[16'h5A25] = 8'hA6;
mem[16'h5A26] = 8'h70;
mem[16'h5A27] = 8'hDE;
mem[16'h5A28] = 8'h75;
mem[16'h5A29] = 8'h5B;
mem[16'h5A2A] = 8'hA6;
mem[16'h5A2B] = 8'h70;
mem[16'h5A2C] = 8'hBD;
mem[16'h5A2D] = 8'h75;
mem[16'h5A2E] = 8'h5B;
mem[16'h5A2F] = 8'hC9;
mem[16'h5A30] = 8'h1D;
mem[16'h5A31] = 8'hD0;
mem[16'h5A32] = 8'h1A;
mem[16'h5A33] = 8'h20;
mem[16'h5A34] = 8'hCD;
mem[16'h5A35] = 8'h75;
mem[16'h5A36] = 8'hA6;
mem[16'h5A37] = 8'h70;
mem[16'h5A38] = 8'hBD;
mem[16'h5A39] = 8'h2C;
mem[16'h5A3A] = 8'h5F;
mem[16'h5A3B] = 8'hC9;
mem[16'h5A3C] = 8'h02;
mem[16'h5A3D] = 8'h90;
mem[16'h5A3E] = 8'hCC;
mem[16'h5A3F] = 8'h38;
mem[16'h5A40] = 8'hE9;
mem[16'h5A41] = 8'h02;
mem[16'h5A42] = 8'h9D;
mem[16'h5A43] = 8'h2C;
mem[16'h5A44] = 8'h5F;
mem[16'h5A45] = 8'h20;
mem[16'h5A46] = 8'h11;
mem[16'h5A47] = 8'h76;
mem[16'h5A48] = 8'hA6;
mem[16'h5A49] = 8'h70;
mem[16'h5A4A] = 8'h4C;
mem[16'h5A4B] = 8'hEA;
mem[16'h5A4C] = 8'h59;
mem[16'h5A4D] = 8'h90;
mem[16'h5A4E] = 8'h15;
mem[16'h5A4F] = 8'hBD;
mem[16'h5A50] = 8'h2C;
mem[16'h5A51] = 8'h5F;
mem[16'h5A52] = 8'hC9;
mem[16'h5A53] = 8'h02;
mem[16'h5A54] = 8'h90;
mem[16'h5A55] = 8'hB5;
mem[16'h5A56] = 8'h38;
mem[16'h5A57] = 8'hE9;
mem[16'h5A58] = 8'h02;
mem[16'h5A59] = 8'h9D;
mem[16'h5A5A] = 8'h2C;
mem[16'h5A5B] = 8'h5F;
mem[16'h5A5C] = 8'h20;
mem[16'h5A5D] = 8'hEB;
mem[16'h5A5E] = 8'h75;
mem[16'h5A5F] = 8'hA6;
mem[16'h5A60] = 8'h70;
mem[16'h5A61] = 8'h4C;
mem[16'h5A62] = 8'hEA;
mem[16'h5A63] = 8'h59;
mem[16'h5A64] = 8'hC9;
mem[16'h5A65] = 8'h16;
mem[16'h5A66] = 8'hB0;
mem[16'h5A67] = 8'hCE;
mem[16'h5A68] = 8'hC9;
mem[16'h5A69] = 8'h15;
mem[16'h5A6A] = 8'hD0;
mem[16'h5A6B] = 8'h15;
mem[16'h5A6C] = 8'h20;
mem[16'h5A6D] = 8'hDC;
mem[16'h5A6E] = 8'h75;
mem[16'h5A6F] = 8'hA6;
mem[16'h5A70] = 8'h70;
mem[16'h5A71] = 8'hBD;
mem[16'h5A72] = 8'h2C;
mem[16'h5A73] = 8'h5F;
mem[16'h5A74] = 8'hC9;
mem[16'h5A75] = 8'h02;
mem[16'h5A76] = 8'h90;
mem[16'h5A77] = 8'h93;
mem[16'h5A78] = 8'h38;
mem[16'h5A79] = 8'hE9;
mem[16'h5A7A] = 8'h02;
mem[16'h5A7B] = 8'h9D;
mem[16'h5A7C] = 8'h2C;
mem[16'h5A7D] = 8'h5F;
mem[16'h5A7E] = 8'h4C;
mem[16'h5A7F] = 8'hEA;
mem[16'h5A80] = 8'h59;
mem[16'h5A81] = 8'hC9;
mem[16'h5A82] = 8'h0F;
mem[16'h5A83] = 8'hB0;
mem[16'h5A84] = 8'hEA;
mem[16'h5A85] = 8'hC9;
mem[16'h5A86] = 8'h0E;
mem[16'h5A87] = 8'hD0;
mem[16'h5A88] = 8'h06;
mem[16'h5A89] = 8'h20;
mem[16'h5A8A] = 8'hDC;
mem[16'h5A8B] = 8'h75;
mem[16'h5A8C] = 8'h4C;
mem[16'h5A8D] = 8'h36;
mem[16'h5A8E] = 8'h5A;
mem[16'h5A8F] = 8'hC9;
mem[16'h5A90] = 8'h08;
mem[16'h5A91] = 8'hB0;
mem[16'h5A92] = 8'hA3;
mem[16'h5A93] = 8'hC9;
mem[16'h5A94] = 8'h07;
mem[16'h5A95] = 8'hF0;
mem[16'h5A96] = 8'h11;
mem[16'h5A97] = 8'hC9;
mem[16'h5A98] = 8'h00;
mem[16'h5A99] = 8'hD0;
mem[16'h5A9A] = 8'hB4;
mem[16'h5A9B] = 8'h20;
mem[16'h5A9C] = 8'hB1;
mem[16'h5A9D] = 8'h75;
mem[16'h5A9E] = 8'hA6;
mem[16'h5A9F] = 8'h70;
mem[16'h5AA0] = 8'hA9;
mem[16'h5AA1] = 8'h00;
mem[16'h5AA2] = 8'h9D;
mem[16'h5AA3] = 8'h75;
mem[16'h5AA4] = 8'h5B;
mem[16'h5AA5] = 8'h4C;
mem[16'h5AA6] = 8'hF6;
mem[16'h5AA7] = 8'h59;
mem[16'h5AA8] = 8'h20;
mem[16'h5AA9] = 8'hCD;
mem[16'h5AAA] = 8'h75;
mem[16'h5AAB] = 8'hA6;
mem[16'h5AAC] = 8'h70;
mem[16'h5AAD] = 8'h4C;
mem[16'h5AAE] = 8'h4F;
mem[16'h5AAF] = 8'h5A;
mem[16'h5AB0] = 8'hAE;
mem[16'h5AB1] = 8'hAF;
mem[16'h5AB2] = 8'h4A;
mem[16'h5AB3] = 8'hCA;
mem[16'h5AB4] = 8'h30;
mem[16'h5AB5] = 8'h2E;
mem[16'h5AB6] = 8'h86;
mem[16'h5AB7] = 8'h70;
mem[16'h5AB8] = 8'hBD;
mem[16'h5AB9] = 8'h75;
mem[16'h5ABA] = 8'h5B;
mem[16'h5ABB] = 8'hD0;
mem[16'h5ABC] = 8'h28;
mem[16'h5ABD] = 8'hBD;
mem[16'h5ABE] = 8'h2C;
mem[16'h5ABF] = 8'h5F;
mem[16'h5AC0] = 8'hC9;
mem[16'h5AC1] = 8'h02;
mem[16'h5AC2] = 8'h90;
mem[16'h5AC3] = 8'h0E;
mem[16'h5AC4] = 8'h38;
mem[16'h5AC5] = 8'hE9;
mem[16'h5AC6] = 8'h02;
mem[16'h5AC7] = 8'h9D;
mem[16'h5AC8] = 8'h2C;
mem[16'h5AC9] = 8'h5F;
mem[16'h5ACA] = 8'h20;
mem[16'h5ACB] = 8'h91;
mem[16'h5ACC] = 8'h5B;
mem[16'h5ACD] = 8'hA6;
mem[16'h5ACE] = 8'h70;
mem[16'h5ACF] = 8'h4C;
mem[16'h5AD0] = 8'hB3;
mem[16'h5AD1] = 8'h5A;
mem[16'h5AD2] = 8'h20;
mem[16'h5AD3] = 8'hC4;
mem[16'h5AD4] = 8'h72;
mem[16'h5AD5] = 8'hA6;
mem[16'h5AD6] = 8'h70;
mem[16'h5AD7] = 8'hA9;
mem[16'h5AD8] = 8'hEB;
mem[16'h5AD9] = 8'h9D;
mem[16'h5ADA] = 8'h2C;
mem[16'h5ADB] = 8'h5F;
mem[16'h5ADC] = 8'h20;
mem[16'h5ADD] = 8'hC4;
mem[16'h5ADE] = 8'h72;
mem[16'h5ADF] = 8'hA6;
mem[16'h5AE0] = 8'h70;
mem[16'h5AE1] = 8'h4C;
mem[16'h5AE2] = 8'hB3;
mem[16'h5AE3] = 8'h5A;
mem[16'h5AE4] = 8'h60;
mem[16'h5AE5] = 8'hC9;
mem[16'h5AE6] = 8'h24;
mem[16'h5AE7] = 8'hD0;
mem[16'h5AE8] = 8'h05;
mem[16'h5AE9] = 8'h20;
mem[16'h5AEA] = 8'hB1;
mem[16'h5AEB] = 8'h75;
mem[16'h5AEC] = 8'hA6;
mem[16'h5AED] = 8'h70;
mem[16'h5AEE] = 8'hDE;
mem[16'h5AEF] = 8'h75;
mem[16'h5AF0] = 8'h5B;
mem[16'h5AF1] = 8'hBD;
mem[16'h5AF2] = 8'h75;
mem[16'h5AF3] = 8'h5B;
mem[16'h5AF4] = 8'hC9;
mem[16'h5AF5] = 8'h1D;
mem[16'h5AF6] = 8'hD0;
mem[16'h5AF7] = 8'h1A;
mem[16'h5AF8] = 8'h20;
mem[16'h5AF9] = 8'hCD;
mem[16'h5AFA] = 8'h75;
mem[16'h5AFB] = 8'hA6;
mem[16'h5AFC] = 8'h70;
mem[16'h5AFD] = 8'hBD;
mem[16'h5AFE] = 8'h2C;
mem[16'h5AFF] = 8'h5F;
mem[16'h5B00] = 8'hC9;
mem[16'h5B01] = 8'h02;
mem[16'h5B02] = 8'h90;
mem[16'h5B03] = 8'hCE;
mem[16'h5B04] = 8'h38;
mem[16'h5B05] = 8'hE9;
mem[16'h5B06] = 8'h02;
mem[16'h5B07] = 8'h9D;
mem[16'h5B08] = 8'h2C;
mem[16'h5B09] = 8'h5F;
mem[16'h5B0A] = 8'h20;
mem[16'h5B0B] = 8'h11;
mem[16'h5B0C] = 8'h76;
mem[16'h5B0D] = 8'hA6;
mem[16'h5B0E] = 8'h70;
mem[16'h5B0F] = 8'h4C;
mem[16'h5B10] = 8'hB3;
mem[16'h5B11] = 8'h5A;
mem[16'h5B12] = 8'h90;
mem[16'h5B13] = 8'h15;
mem[16'h5B14] = 8'hBD;
mem[16'h5B15] = 8'h2C;
mem[16'h5B16] = 8'h5F;
mem[16'h5B17] = 8'hC9;
mem[16'h5B18] = 8'h02;
mem[16'h5B19] = 8'h90;
mem[16'h5B1A] = 8'hB7;
mem[16'h5B1B] = 8'h38;
mem[16'h5B1C] = 8'hE9;
mem[16'h5B1D] = 8'h02;
mem[16'h5B1E] = 8'h9D;
mem[16'h5B1F] = 8'h2C;
mem[16'h5B20] = 8'h5F;
mem[16'h5B21] = 8'h20;
mem[16'h5B22] = 8'hEB;
mem[16'h5B23] = 8'h75;
mem[16'h5B24] = 8'hA6;
mem[16'h5B25] = 8'h70;
mem[16'h5B26] = 8'h4C;
mem[16'h5B27] = 8'hB3;
mem[16'h5B28] = 8'h5A;
mem[16'h5B29] = 8'hC9;
mem[16'h5B2A] = 8'h16;
mem[16'h5B2B] = 8'hB0;
mem[16'h5B2C] = 8'hCE;
mem[16'h5B2D] = 8'hC9;
mem[16'h5B2E] = 8'h15;
mem[16'h5B2F] = 8'hD0;
mem[16'h5B30] = 8'h15;
mem[16'h5B31] = 8'h20;
mem[16'h5B32] = 8'hDC;
mem[16'h5B33] = 8'h75;
mem[16'h5B34] = 8'hA6;
mem[16'h5B35] = 8'h70;
mem[16'h5B36] = 8'hBD;
mem[16'h5B37] = 8'h2C;
mem[16'h5B38] = 8'h5F;
mem[16'h5B39] = 8'hC9;
mem[16'h5B3A] = 8'h02;
mem[16'h5B3B] = 8'h90;
mem[16'h5B3C] = 8'h95;
mem[16'h5B3D] = 8'h38;
mem[16'h5B3E] = 8'hE9;
mem[16'h5B3F] = 8'h02;
mem[16'h5B40] = 8'h9D;
mem[16'h5B41] = 8'h2C;
mem[16'h5B42] = 8'h5F;
mem[16'h5B43] = 8'h4C;
mem[16'h5B44] = 8'hB3;
mem[16'h5B45] = 8'h5A;
mem[16'h5B46] = 8'hC9;
mem[16'h5B47] = 8'h0F;
mem[16'h5B48] = 8'hB0;
mem[16'h5B49] = 8'hEA;
mem[16'h5B4A] = 8'hC9;
mem[16'h5B4B] = 8'h0E;
mem[16'h5B4C] = 8'hD0;
mem[16'h5B4D] = 8'h06;
mem[16'h5B4E] = 8'h20;
mem[16'h5B4F] = 8'hDC;
mem[16'h5B50] = 8'h75;
mem[16'h5B51] = 8'h4C;
mem[16'h5B52] = 8'hFB;
mem[16'h5B53] = 8'h5A;
mem[16'h5B54] = 8'hC9;
mem[16'h5B55] = 8'h08;
mem[16'h5B56] = 8'hB0;
mem[16'h5B57] = 8'hA3;
mem[16'h5B58] = 8'hC9;
mem[16'h5B59] = 8'h07;
mem[16'h5B5A] = 8'hF0;
mem[16'h5B5B] = 8'h11;
mem[16'h5B5C] = 8'hC9;
mem[16'h5B5D] = 8'h00;
mem[16'h5B5E] = 8'hD0;
mem[16'h5B5F] = 8'hB4;
mem[16'h5B60] = 8'h20;
mem[16'h5B61] = 8'hB1;
mem[16'h5B62] = 8'h75;
mem[16'h5B63] = 8'hA6;
mem[16'h5B64] = 8'h70;
mem[16'h5B65] = 8'hA9;
mem[16'h5B66] = 8'h00;
mem[16'h5B67] = 8'h9D;
mem[16'h5B68] = 8'h75;
mem[16'h5B69] = 8'h5B;
mem[16'h5B6A] = 8'h4C;
mem[16'h5B6B] = 8'hBD;
mem[16'h5B6C] = 8'h5A;
mem[16'h5B6D] = 8'h20;
mem[16'h5B6E] = 8'hCD;
mem[16'h5B6F] = 8'h75;
mem[16'h5B70] = 8'hA6;
mem[16'h5B71] = 8'h70;
mem[16'h5B72] = 8'h4C;
mem[16'h5B73] = 8'h14;
mem[16'h5B74] = 8'h5B;
mem[16'h5B75] = 8'h00;
mem[16'h5B76] = 8'h00;
mem[16'h5B77] = 8'h00;
mem[16'h5B78] = 8'h00;
mem[16'h5B79] = 8'h00;
mem[16'h5B7A] = 8'h00;
mem[16'h5B7B] = 8'h00;
mem[16'h5B7C] = 8'h00;
mem[16'h5B7D] = 8'h00;
mem[16'h5B7E] = 8'h00;
mem[16'h5B7F] = 8'h00;
mem[16'h5B80] = 8'h00;
mem[16'h5B81] = 8'h00;
mem[16'h5B82] = 8'h00;
mem[16'h5B83] = 8'h07;
mem[16'h5B84] = 8'h07;
mem[16'h5B85] = 8'h07;
mem[16'h5B86] = 8'h07;
mem[16'h5B87] = 8'h07;
mem[16'h5B88] = 8'h07;
mem[16'h5B89] = 8'h07;
mem[16'h5B8A] = 8'h07;
mem[16'h5B8B] = 8'h07;
mem[16'h5B8C] = 8'h07;
mem[16'h5B8D] = 8'h07;
mem[16'h5B8E] = 8'h07;
mem[16'h5B8F] = 8'h07;
mem[16'h5B90] = 8'h07;
mem[16'h5B91] = 8'hA6;
mem[16'h5B92] = 8'h70;
mem[16'h5B93] = 8'hBD;
mem[16'h5B94] = 8'h1E;
mem[16'h5B95] = 8'h5F;
mem[16'h5B96] = 8'h85;
mem[16'h5B97] = 8'h56;
mem[16'h5B98] = 8'hBC;
mem[16'h5B99] = 8'h2C;
mem[16'h5B9A] = 8'h5F;
mem[16'h5B9B] = 8'h84;
mem[16'h5B9C] = 8'h57;
mem[16'h5B9D] = 8'hB9;
mem[16'h5B9E] = 8'h3E;
mem[16'h5B9F] = 8'h8C;
mem[16'h5BA0] = 8'hAA;
mem[16'h5BA1] = 8'hBD;
mem[16'h5BA2] = 8'h94;
mem[16'h5BA3] = 8'h8E;
mem[16'h5BA4] = 8'hAA;
mem[16'h5BA5] = 8'hA4;
mem[16'h5BA6] = 8'h70;
mem[16'h5BA7] = 8'hB9;
mem[16'h5BA8] = 8'h83;
mem[16'h5BA9] = 8'h5B;
mem[16'h5BAA] = 8'hF0;
mem[16'h5BAB] = 8'h29;
mem[16'h5BAC] = 8'hC9;
mem[16'h5BAD] = 8'h08;
mem[16'h5BAE] = 8'hF0;
mem[16'h5BAF] = 8'h37;
mem[16'h5BB0] = 8'h90;
mem[16'h5BB1] = 8'h2C;
mem[16'h5BB2] = 8'hBD;
mem[16'h5BB3] = 8'h0C;
mem[16'h5BB4] = 8'h5C;
mem[16'h5BB5] = 8'hBC;
mem[16'h5BB6] = 8'h13;
mem[16'h5BB7] = 8'h5C;
mem[16'h5BB8] = 8'h20;
mem[16'h5BB9] = 8'hD1;
mem[16'h5BBA] = 8'h8A;
mem[16'h5BBB] = 8'hA9;
mem[16'h5BBC] = 8'h2C;
mem[16'h5BBD] = 8'h8D;
mem[16'h5BBE] = 8'hCA;
mem[16'h5BBF] = 8'h8A;
mem[16'h5BC0] = 8'h20;
mem[16'h5BC1] = 8'h79;
mem[16'h5BC2] = 8'h8A;
mem[16'h5BC3] = 8'hA6;
mem[16'h5BC4] = 8'h70;
mem[16'h5BC5] = 8'hFE;
mem[16'h5BC6] = 8'h83;
mem[16'h5BC7] = 8'h5B;
mem[16'h5BC8] = 8'hBD;
mem[16'h5BC9] = 8'h83;
mem[16'h5BCA] = 8'h5B;
mem[16'h5BCB] = 8'hC9;
mem[16'h5BCC] = 8'h18;
mem[16'h5BCD] = 8'h90;
mem[16'h5BCE] = 8'h05;
mem[16'h5BCF] = 8'hA9;
mem[16'h5BD0] = 8'h00;
mem[16'h5BD1] = 8'h9D;
mem[16'h5BD2] = 8'h83;
mem[16'h5BD3] = 8'h5B;
mem[16'h5BD4] = 8'h60;
mem[16'h5BD5] = 8'hBD;
mem[16'h5BD6] = 8'hF0;
mem[16'h5BD7] = 8'h5B;
mem[16'h5BD8] = 8'hBC;
mem[16'h5BD9] = 8'hF7;
mem[16'h5BDA] = 8'h5B;
mem[16'h5BDB] = 8'h4C;
mem[16'h5BDC] = 8'hB8;
mem[16'h5BDD] = 8'h5B;
mem[16'h5BDE] = 8'hBD;
mem[16'h5BDF] = 8'hFE;
mem[16'h5BE0] = 8'h5B;
mem[16'h5BE1] = 8'hBC;
mem[16'h5BE2] = 8'h05;
mem[16'h5BE3] = 8'h5C;
mem[16'h5BE4] = 8'h4C;
mem[16'h5BE5] = 8'hB8;
mem[16'h5BE6] = 8'h5B;
mem[16'h5BE7] = 8'hBD;
mem[16'h5BE8] = 8'h1A;
mem[16'h5BE9] = 8'h5C;
mem[16'h5BEA] = 8'hBC;
mem[16'h5BEB] = 8'h21;
mem[16'h5BEC] = 8'h5C;
mem[16'h5BED] = 8'h4C;
mem[16'h5BEE] = 8'hB8;
mem[16'h5BEF] = 8'h5B;
mem[16'h5BF0] = 8'h5E;
mem[16'h5BF1] = 8'h32;
mem[16'h5BF2] = 8'h06;
mem[16'h5BF3] = 8'hDA;
mem[16'h5BF4] = 8'hAE;
mem[16'h5BF5] = 8'h82;
mem[16'h5BF6] = 8'h56;
mem[16'h5BF7] = 8'h7D;
mem[16'h5BF8] = 8'h7D;
mem[16'h5BF9] = 8'h7D;
mem[16'h5BFA] = 8'h7C;
mem[16'h5BFB] = 8'h7C;
mem[16'h5BFC] = 8'h7C;
mem[16'h5BFD] = 8'h7C;
mem[16'h5BFE] = 8'h92;
mem[16'h5BFF] = 8'h66;
mem[16'h5C00] = 8'h3A;
mem[16'h5C01] = 8'h0E;
mem[16'h5C02] = 8'hE2;
mem[16'h5C03] = 8'hB6;
mem[16'h5C04] = 8'h8A;
mem[16'h5C05] = 8'h7E;
mem[16'h5C06] = 8'h7E;
mem[16'h5C07] = 8'h7E;
mem[16'h5C08] = 8'h7E;
mem[16'h5C09] = 8'h7D;
mem[16'h5C0A] = 8'h7D;
mem[16'h5C0B] = 8'h7D;
mem[16'h5C0C] = 8'h32;
mem[16'h5C0D] = 8'h5E;
mem[16'h5C0E] = 8'h8A;
mem[16'h5C0F] = 8'hB6;
mem[16'h5C10] = 8'hE2;
mem[16'h5C11] = 8'h0E;
mem[16'h5C12] = 8'h3A;
mem[16'h5C13] = 8'h61;
mem[16'h5C14] = 8'h61;
mem[16'h5C15] = 8'h61;
mem[16'h5C16] = 8'h61;
mem[16'h5C17] = 8'h61;
mem[16'h5C18] = 8'h62;
mem[16'h5C19] = 8'h62;
mem[16'h5C1A] = 8'hBD;
mem[16'h5C1B] = 8'h91;
mem[16'h5C1C] = 8'h65;
mem[16'h5C1D] = 8'h39;
mem[16'h5C1E] = 8'h0D;
mem[16'h5C1F] = 8'hE1;
mem[16'h5C20] = 8'hB5;
mem[16'h5C21] = 8'h93;
mem[16'h5C22] = 8'h93;
mem[16'h5C23] = 8'h93;
mem[16'h5C24] = 8'h93;
mem[16'h5C25] = 8'h93;
mem[16'h5C26] = 8'h92;
mem[16'h5C27] = 8'h92;
mem[16'h5C28] = 8'hAE;
mem[16'h5C29] = 8'hAD;
mem[16'h5C2A] = 8'h4A;
mem[16'h5C2B] = 8'hCA;
mem[16'h5C2C] = 8'h30;
mem[16'h5C2D] = 8'h33;
mem[16'h5C2E] = 8'h86;
mem[16'h5C2F] = 8'h70;
mem[16'h5C30] = 8'hBC;
mem[16'h5C31] = 8'hAF;
mem[16'h5C32] = 8'h60;
mem[16'h5C33] = 8'h84;
mem[16'h5C34] = 8'h57;
mem[16'h5C35] = 8'hBD;
mem[16'h5C36] = 8'hB3;
mem[16'h5C37] = 8'h60;
mem[16'h5C38] = 8'h85;
mem[16'h5C39] = 8'h56;
mem[16'h5C3A] = 8'h20;
mem[16'h5C3B] = 8'h92;
mem[16'h5C3C] = 8'h5C;
mem[16'h5C3D] = 8'hA6;
mem[16'h5C3E] = 8'h70;
mem[16'h5C3F] = 8'hBD;
mem[16'h5C40] = 8'hAF;
mem[16'h5C41] = 8'h60;
mem[16'h5C42] = 8'h18;
mem[16'h5C43] = 8'h69;
mem[16'h5C44] = 8'h02;
mem[16'h5C45] = 8'h9D;
mem[16'h5C46] = 8'hAF;
mem[16'h5C47] = 8'h60;
mem[16'h5C48] = 8'hC9;
mem[16'h5C49] = 8'hFE;
mem[16'h5C4A] = 8'h90;
mem[16'h5C4B] = 8'hDF;
mem[16'h5C4C] = 8'h20;
mem[16'h5C4D] = 8'h4D;
mem[16'h5C4E] = 8'h60;
mem[16'h5C4F] = 8'hA6;
mem[16'h5C50] = 8'h70;
mem[16'h5C51] = 8'hBD;
mem[16'h5C52] = 8'hB3;
mem[16'h5C53] = 8'h60;
mem[16'h5C54] = 8'h29;
mem[16'h5C55] = 8'h01;
mem[16'h5C56] = 8'h9D;
mem[16'h5C57] = 8'hAF;
mem[16'h5C58] = 8'h60;
mem[16'h5C59] = 8'h20;
mem[16'h5C5A] = 8'h4D;
mem[16'h5C5B] = 8'h60;
mem[16'h5C5C] = 8'hA6;
mem[16'h5C5D] = 8'h70;
mem[16'h5C5E] = 8'h4C;
mem[16'h5C5F] = 8'h2B;
mem[16'h5C60] = 8'h5C;
mem[16'h5C61] = 8'h60;
mem[16'h5C62] = 8'hAE;
mem[16'h5C63] = 8'hAA;
mem[16'h5C64] = 8'h4A;
mem[16'h5C65] = 8'hCA;
mem[16'h5C66] = 8'h30;
mem[16'h5C67] = 8'h29;
mem[16'h5C68] = 8'h86;
mem[16'h5C69] = 8'h70;
mem[16'h5C6A] = 8'h20;
mem[16'h5C6B] = 8'hBA;
mem[16'h5C6C] = 8'h5C;
mem[16'h5C6D] = 8'hA6;
mem[16'h5C6E] = 8'h70;
mem[16'h5C6F] = 8'hBD;
mem[16'h5C70] = 8'hA7;
mem[16'h5C71] = 8'h60;
mem[16'h5C72] = 8'h18;
mem[16'h5C73] = 8'h69;
mem[16'h5C74] = 8'h02;
mem[16'h5C75] = 8'h9D;
mem[16'h5C76] = 8'hA7;
mem[16'h5C77] = 8'h60;
mem[16'h5C78] = 8'hC9;
mem[16'h5C79] = 8'hFE;
mem[16'h5C7A] = 8'h90;
mem[16'h5C7B] = 8'hE9;
mem[16'h5C7C] = 8'h20;
mem[16'h5C7D] = 8'h69;
mem[16'h5C7E] = 8'h60;
mem[16'h5C7F] = 8'hA6;
mem[16'h5C80] = 8'h70;
mem[16'h5C81] = 8'hBD;
mem[16'h5C82] = 8'hAB;
mem[16'h5C83] = 8'h60;
mem[16'h5C84] = 8'h29;
mem[16'h5C85] = 8'h01;
mem[16'h5C86] = 8'h9D;
mem[16'h5C87] = 8'hA7;
mem[16'h5C88] = 8'h60;
mem[16'h5C89] = 8'h20;
mem[16'h5C8A] = 8'h69;
mem[16'h5C8B] = 8'h60;
mem[16'h5C8C] = 8'hA6;
mem[16'h5C8D] = 8'h70;
mem[16'h5C8E] = 8'h4C;
mem[16'h5C8F] = 8'h65;
mem[16'h5C90] = 8'h5C;
mem[16'h5C91] = 8'h60;
mem[16'h5C92] = 8'hB9;
mem[16'h5C93] = 8'h3E;
mem[16'h5C94] = 8'h8C;
mem[16'h5C95] = 8'hAA;
mem[16'h5C96] = 8'hBD;
mem[16'h5C97] = 8'h94;
mem[16'h5C98] = 8'h8E;
mem[16'h5C99] = 8'hAA;
mem[16'h5C9A] = 8'hBD;
mem[16'h5C9B] = 8'hAC;
mem[16'h5C9C] = 8'h5C;
mem[16'h5C9D] = 8'hBC;
mem[16'h5C9E] = 8'hB3;
mem[16'h5C9F] = 8'h5C;
mem[16'h5CA0] = 8'h20;
mem[16'h5CA1] = 8'h3B;
mem[16'h5CA2] = 8'h8B;
mem[16'h5CA3] = 8'hA9;
mem[16'h5CA4] = 8'h18;
mem[16'h5CA5] = 8'h8D;
mem[16'h5CA6] = 8'h34;
mem[16'h5CA7] = 8'h8B;
mem[16'h5CA8] = 8'h20;
mem[16'h5CA9] = 8'hF0;
mem[16'h5CAA] = 8'h8A;
mem[16'h5CAB] = 8'h60;
mem[16'h5CAC] = 8'hEE;
mem[16'h5CAD] = 8'h06;
mem[16'h5CAE] = 8'h1E;
mem[16'h5CAF] = 8'h36;
mem[16'h5CB0] = 8'h4E;
mem[16'h5CB1] = 8'h66;
mem[16'h5CB2] = 8'h7E;
mem[16'h5CB3] = 8'h5C;
mem[16'h5CB4] = 8'h5D;
mem[16'h5CB5] = 8'h5D;
mem[16'h5CB6] = 8'h5D;
mem[16'h5CB7] = 8'h5D;
mem[16'h5CB8] = 8'h5D;
mem[16'h5CB9] = 8'h5D;
mem[16'h5CBA] = 8'hA6;
mem[16'h5CBB] = 8'h70;
mem[16'h5CBC] = 8'hBD;
mem[16'h5CBD] = 8'hAB;
mem[16'h5CBE] = 8'h60;
mem[16'h5CBF] = 8'h85;
mem[16'h5CC0] = 8'h56;
mem[16'h5CC1] = 8'hBC;
mem[16'h5CC2] = 8'hA7;
mem[16'h5CC3] = 8'h60;
mem[16'h5CC4] = 8'h84;
mem[16'h5CC5] = 8'h57;
mem[16'h5CC6] = 8'hB9;
mem[16'h5CC7] = 8'h3E;
mem[16'h5CC8] = 8'h8C;
mem[16'h5CC9] = 8'hAA;
mem[16'h5CCA] = 8'hBD;
mem[16'h5CCB] = 8'h94;
mem[16'h5CCC] = 8'h8E;
mem[16'h5CCD] = 8'hAA;
mem[16'h5CCE] = 8'hBD;
mem[16'h5CCF] = 8'hE0;
mem[16'h5CD0] = 8'h5C;
mem[16'h5CD1] = 8'hBC;
mem[16'h5CD2] = 8'hE7;
mem[16'h5CD3] = 8'h5C;
mem[16'h5CD4] = 8'h20;
mem[16'h5CD5] = 8'h3B;
mem[16'h5CD6] = 8'h8B;
mem[16'h5CD7] = 8'hA9;
mem[16'h5CD8] = 8'h1B;
mem[16'h5CD9] = 8'h8D;
mem[16'h5CDA] = 8'h34;
mem[16'h5CDB] = 8'h8B;
mem[16'h5CDC] = 8'h20;
mem[16'h5CDD] = 8'hF0;
mem[16'h5CDE] = 8'h8A;
mem[16'h5CDF] = 8'h60;
mem[16'h5CE0] = 8'hA9;
mem[16'h5CE1] = 8'h8E;
mem[16'h5CE2] = 8'h73;
mem[16'h5CE3] = 8'h58;
mem[16'h5CE4] = 8'h3D;
mem[16'h5CE5] = 8'h22;
mem[16'h5CE6] = 8'h07;
mem[16'h5CE7] = 8'h72;
mem[16'h5CE8] = 8'h72;
mem[16'h5CE9] = 8'h72;
mem[16'h5CEA] = 8'h72;
mem[16'h5CEB] = 8'h72;
mem[16'h5CEC] = 8'h72;
mem[16'h5CED] = 8'h72;
mem[16'h5CEE] = 8'hB6;
mem[16'h5CEF] = 8'h58;
mem[16'h5CF0] = 8'h01;
mem[16'h5CF1] = 8'hB6;
mem[16'h5CF2] = 8'h58;
mem[16'h5CF3] = 8'h01;
mem[16'h5CF4] = 8'hD4;
mem[16'h5CF5] = 8'h58;
mem[16'h5CF6] = 8'h00;
mem[16'h5CF7] = 8'h84;
mem[16'h5CF8] = 8'h00;
mem[16'h5CF9] = 8'h01;
mem[16'h5CFA] = 8'h8B;
mem[16'h5CFB] = 8'h00;
mem[16'h5CFC] = 8'h01;
mem[16'h5CFD] = 8'hD4;
mem[16'h5CFE] = 8'h58;
mem[16'h5CFF] = 8'h00;
mem[16'h5D00] = 8'hB6;
mem[16'h5D01] = 8'h58;
mem[16'h5D02] = 8'h01;
mem[16'h5D03] = 8'hB6;
mem[16'h5D04] = 8'h58;
mem[16'h5D05] = 8'h01;
mem[16'h5D06] = 8'hEC;
mem[16'h5D07] = 8'h30;
mem[16'h5D08] = 8'h03;
mem[16'h5D09] = 8'hEC;
mem[16'h5D0A] = 8'h30;
mem[16'h5D0B] = 8'h03;
mem[16'h5D0C] = 8'hA8;
mem[16'h5D0D] = 8'h31;
mem[16'h5D0E] = 8'h01;
mem[16'h5D0F] = 8'h88;
mem[16'h5D10] = 8'h00;
mem[16'h5D11] = 8'h02;
mem[16'h5D12] = 8'h96;
mem[16'h5D13] = 8'h00;
mem[16'h5D14] = 8'h02;
mem[16'h5D15] = 8'hA8;
mem[16'h5D16] = 8'h31;
mem[16'h5D17] = 8'h01;
mem[16'h5D18] = 8'hEC;
mem[16'h5D19] = 8'h30;
mem[16'h5D1A] = 8'h03;
mem[16'h5D1B] = 8'hEC;
mem[16'h5D1C] = 8'h30;
mem[16'h5D1D] = 8'h03;
mem[16'h5D1E] = 8'hD8;
mem[16'h5D1F] = 8'h61;
mem[16'h5D20] = 8'h06;
mem[16'h5D21] = 8'hD8;
mem[16'h5D22] = 8'h61;
mem[16'h5D23] = 8'h06;
mem[16'h5D24] = 8'hD0;
mem[16'h5D25] = 8'h62;
mem[16'h5D26] = 8'h02;
mem[16'h5D27] = 8'h90;
mem[16'h5D28] = 8'h00;
mem[16'h5D29] = 8'h04;
mem[16'h5D2A] = 8'hAC;
mem[16'h5D2B] = 8'h00;
mem[16'h5D2C] = 8'h04;
mem[16'h5D2D] = 8'hD0;
mem[16'h5D2E] = 8'h62;
mem[16'h5D2F] = 8'h02;
mem[16'h5D30] = 8'hD8;
mem[16'h5D31] = 8'h61;
mem[16'h5D32] = 8'h06;
mem[16'h5D33] = 8'hD8;
mem[16'h5D34] = 8'h61;
mem[16'h5D35] = 8'h06;
mem[16'h5D36] = 8'hB0;
mem[16'h5D37] = 8'h43;
mem[16'h5D38] = 8'h0D;
mem[16'h5D39] = 8'hB0;
mem[16'h5D3A] = 8'h43;
mem[16'h5D3B] = 8'h0D;
mem[16'h5D3C] = 8'hA0;
mem[16'h5D3D] = 8'h45;
mem[16'h5D3E] = 8'h05;
mem[16'h5D3F] = 8'hA0;
mem[16'h5D40] = 8'h00;
mem[16'h5D41] = 8'h08;
mem[16'h5D42] = 8'hD8;
mem[16'h5D43] = 8'h00;
mem[16'h5D44] = 8'h08;
mem[16'h5D45] = 8'hA0;
mem[16'h5D46] = 8'h45;
mem[16'h5D47] = 8'h05;
mem[16'h5D48] = 8'hB0;
mem[16'h5D49] = 8'h43;
mem[16'h5D4A] = 8'h0D;
mem[16'h5D4B] = 8'hB0;
mem[16'h5D4C] = 8'h43;
mem[16'h5D4D] = 8'h0D;
mem[16'h5D4E] = 8'hE0;
mem[16'h5D4F] = 8'h06;
mem[16'h5D50] = 8'h1B;
mem[16'h5D51] = 8'hE0;
mem[16'h5D52] = 8'h06;
mem[16'h5D53] = 8'h1B;
mem[16'h5D54] = 8'hC0;
mem[16'h5D55] = 8'h0A;
mem[16'h5D56] = 8'h0B;
mem[16'h5D57] = 8'hC0;
mem[16'h5D58] = 8'h00;
mem[16'h5D59] = 8'h10;
mem[16'h5D5A] = 8'hB0;
mem[16'h5D5B] = 8'h01;
mem[16'h5D5C] = 8'h10;
mem[16'h5D5D] = 8'hC0;
mem[16'h5D5E] = 8'h0A;
mem[16'h5D5F] = 8'h0B;
mem[16'h5D60] = 8'hE0;
mem[16'h5D61] = 8'h06;
mem[16'h5D62] = 8'h1B;
mem[16'h5D63] = 8'hE0;
mem[16'h5D64] = 8'h06;
mem[16'h5D65] = 8'h1B;
mem[16'h5D66] = 8'hC0;
mem[16'h5D67] = 8'h0D;
mem[16'h5D68] = 8'h36;
mem[16'h5D69] = 8'hC0;
mem[16'h5D6A] = 8'h0D;
mem[16'h5D6B] = 8'h36;
mem[16'h5D6C] = 8'h80;
mem[16'h5D6D] = 8'h15;
mem[16'h5D6E] = 8'h16;
mem[16'h5D6F] = 8'h80;
mem[16'h5D70] = 8'h01;
mem[16'h5D71] = 8'h20;
mem[16'h5D72] = 8'hE0;
mem[16'h5D73] = 8'h02;
mem[16'h5D74] = 8'h20;
mem[16'h5D75] = 8'h80;
mem[16'h5D76] = 8'h15;
mem[16'h5D77] = 8'h16;
mem[16'h5D78] = 8'hC0;
mem[16'h5D79] = 8'h0D;
mem[16'h5D7A] = 8'h36;
mem[16'h5D7B] = 8'hC0;
mem[16'h5D7C] = 8'h0D;
mem[16'h5D7D] = 8'h36;
mem[16'h5D7E] = 8'h80;
mem[16'h5D7F] = 8'h1B;
mem[16'h5D80] = 8'h6C;
mem[16'h5D81] = 8'h80;
mem[16'h5D82] = 8'h1B;
mem[16'h5D83] = 8'h6C;
mem[16'h5D84] = 8'h80;
mem[16'h5D85] = 8'h2A;
mem[16'h5D86] = 8'h2C;
mem[16'h5D87] = 8'h80;
mem[16'h5D88] = 8'h02;
mem[16'h5D89] = 8'h40;
mem[16'h5D8A] = 8'hC0;
mem[16'h5D8B] = 8'h05;
mem[16'h5D8C] = 8'h40;
mem[16'h5D8D] = 8'h80;
mem[16'h5D8E] = 8'h2A;
mem[16'h5D8F] = 8'h2C;
mem[16'h5D90] = 8'h80;
mem[16'h5D91] = 8'h1B;
mem[16'h5D92] = 8'h6C;
mem[16'h5D93] = 8'h80;
mem[16'h5D94] = 8'h1B;
mem[16'h5D95] = 8'h6C;
mem[16'h5D96] = 8'h20;
mem[16'h5D97] = 8'h9C;
mem[16'h5D98] = 8'h5F;
mem[16'h5D99] = 8'h20;
mem[16'h5D9A] = 8'hD7;
mem[16'h5D9B] = 8'h5D;
mem[16'h5D9C] = 8'h20;
mem[16'h5D9D] = 8'h6B;
mem[16'h5D9E] = 8'h5F;
mem[16'h5D9F] = 8'h20;
mem[16'h5DA0] = 8'h3A;
mem[16'h5DA1] = 8'h5F;
mem[16'h5DA2] = 8'h20;
mem[16'h5DA3] = 8'hA6;
mem[16'h5DA4] = 8'h5D;
mem[16'h5DA5] = 8'h60;
mem[16'h5DA6] = 8'hAE;
mem[16'h5DA7] = 8'hAE;
mem[16'h5DA8] = 8'h4A;
mem[16'h5DA9] = 8'h8A;
mem[16'h5DAA] = 8'h38;
mem[16'h5DAB] = 8'hE9;
mem[16'h5DAC] = 8'h01;
mem[16'h5DAD] = 8'h85;
mem[16'h5DAE] = 8'h6E;
mem[16'h5DAF] = 8'hCA;
mem[16'h5DB0] = 8'h30;
mem[16'h5DB1] = 8'h24;
mem[16'h5DB2] = 8'h86;
mem[16'h5DB3] = 8'h70;
mem[16'h5DB4] = 8'hA9;
mem[16'h5DB5] = 8'h6C;
mem[16'h5DB6] = 8'h9D;
mem[16'h5DB7] = 8'h4A;
mem[16'h5DB8] = 8'h60;
mem[16'h5DB9] = 8'hE4;
mem[16'h5DBA] = 8'h6E;
mem[16'h5DBB] = 8'h90;
mem[16'h5DBC] = 8'h08;
mem[16'h5DBD] = 8'hA9;
mem[16'h5DBE] = 8'h0E;
mem[16'h5DBF] = 8'h9D;
mem[16'h5DC0] = 8'h47;
mem[16'h5DC1] = 8'h60;
mem[16'h5DC2] = 8'h4C;
mem[16'h5DC3] = 8'hCE;
mem[16'h5DC4] = 8'h5D;
mem[16'h5DC5] = 8'hBD;
mem[16'h5DC6] = 8'h48;
mem[16'h5DC7] = 8'h60;
mem[16'h5DC8] = 8'h18;
mem[16'h5DC9] = 8'h69;
mem[16'h5DCA] = 8'h62;
mem[16'h5DCB] = 8'h9D;
mem[16'h5DCC] = 8'h47;
mem[16'h5DCD] = 8'h60;
mem[16'h5DCE] = 8'h20;
mem[16'h5DCF] = 8'h13;
mem[16'h5DD0] = 8'h60;
mem[16'h5DD1] = 8'hA6;
mem[16'h5DD2] = 8'h70;
mem[16'h5DD3] = 8'h4C;
mem[16'h5DD4] = 8'hAF;
mem[16'h5DD5] = 8'h5D;
mem[16'h5DD6] = 8'h60;
mem[16'h5DD7] = 8'hAE;
mem[16'h5DD8] = 8'hAB;
mem[16'h5DD9] = 8'h4A;
mem[16'h5DDA] = 8'hCA;
mem[16'h5DDB] = 8'h30;
mem[16'h5DDC] = 8'h27;
mem[16'h5DDD] = 8'h86;
mem[16'h5DDE] = 8'h70;
mem[16'h5DDF] = 8'hA9;
mem[16'h5DE0] = 8'h87;
mem[16'h5DE1] = 8'h9D;
mem[16'h5DE2] = 8'hEF;
mem[16'h5DE3] = 8'h60;
mem[16'h5DE4] = 8'hE8;
mem[16'h5DE5] = 8'hEC;
mem[16'h5DE6] = 8'hAB;
mem[16'h5DE7] = 8'h4A;
mem[16'h5DE8] = 8'hCA;
mem[16'h5DE9] = 8'h90;
mem[16'h5DEA] = 8'h08;
mem[16'h5DEB] = 8'hA9;
mem[16'h5DEC] = 8'h23;
mem[16'h5DED] = 8'h9D;
mem[16'h5DEE] = 8'hEB;
mem[16'h5DEF] = 8'h60;
mem[16'h5DF0] = 8'h4C;
mem[16'h5DF1] = 8'hFC;
mem[16'h5DF2] = 8'h5D;
mem[16'h5DF3] = 8'hBD;
mem[16'h5DF4] = 8'hEC;
mem[16'h5DF5] = 8'h60;
mem[16'h5DF6] = 8'h18;
mem[16'h5DF7] = 8'h69;
mem[16'h5DF8] = 8'h54;
mem[16'h5DF9] = 8'h9D;
mem[16'h5DFA] = 8'hEB;
mem[16'h5DFB] = 8'h60;
mem[16'h5DFC] = 8'h20;
mem[16'h5DFD] = 8'hB7;
mem[16'h5DFE] = 8'h60;
mem[16'h5DFF] = 8'hA6;
mem[16'h5E00] = 8'h70;
mem[16'h5E01] = 8'h4C;
mem[16'h5E02] = 8'hDA;
mem[16'h5E03] = 8'h5D;
mem[16'h5E04] = 8'h60;
mem[16'h5E05] = 8'hAD;
mem[16'h5E06] = 8'hAF;
mem[16'h5E07] = 8'h4A;
mem[16'h5E08] = 8'hAA;
mem[16'h5E09] = 8'hCA;
mem[16'h5E0A] = 8'hA9;
mem[16'h5E0B] = 8'h25;
mem[16'h5E0C] = 8'h9D;
mem[16'h5E0D] = 8'h1E;
mem[16'h5E0E] = 8'h5F;
mem[16'h5E0F] = 8'hA9;
mem[16'h5E10] = 8'h03;
mem[16'h5E11] = 8'h9D;
mem[16'h5E12] = 8'h2C;
mem[16'h5E13] = 8'h5F;
mem[16'h5E14] = 8'h86;
mem[16'h5E15] = 8'h70;
mem[16'h5E16] = 8'h20;
mem[16'h5E17] = 8'hC6;
mem[16'h5E18] = 8'h5E;
mem[16'h5E19] = 8'hAD;
mem[16'h5E1A] = 8'hAF;
mem[16'h5E1B] = 8'h4A;
mem[16'h5E1C] = 8'hAA;
mem[16'h5E1D] = 8'hCA;
mem[16'h5E1E] = 8'h38;
mem[16'h5E1F] = 8'hED;
mem[16'h5E20] = 8'h63;
mem[16'h5E21] = 8'h5E;
mem[16'h5E22] = 8'h8D;
mem[16'h5E23] = 8'hC5;
mem[16'h5E24] = 8'h5E;
mem[16'h5E25] = 8'hCA;
mem[16'h5E26] = 8'hA9;
mem[16'h5E27] = 8'h25;
mem[16'h5E28] = 8'h9D;
mem[16'h5E29] = 8'h1E;
mem[16'h5E2A] = 8'h5F;
mem[16'h5E2B] = 8'hBD;
mem[16'h5E2C] = 8'h2D;
mem[16'h5E2D] = 8'h5F;
mem[16'h5E2E] = 8'h18;
mem[16'h5E2F] = 8'h69;
mem[16'h5E30] = 8'h12;
mem[16'h5E31] = 8'h9D;
mem[16'h5E32] = 8'h2C;
mem[16'h5E33] = 8'h5F;
mem[16'h5E34] = 8'h86;
mem[16'h5E35] = 8'h70;
mem[16'h5E36] = 8'h20;
mem[16'h5E37] = 8'hC6;
mem[16'h5E38] = 8'h5E;
mem[16'h5E39] = 8'hA6;
mem[16'h5E3A] = 8'h70;
mem[16'h5E3B] = 8'hEC;
mem[16'h5E3C] = 8'hC5;
mem[16'h5E3D] = 8'h5E;
mem[16'h5E3E] = 8'hF0;
mem[16'h5E3F] = 8'h03;
mem[16'h5E40] = 8'h4C;
mem[16'h5E41] = 8'h25;
mem[16'h5E42] = 8'h5E;
mem[16'h5E43] = 8'hCA;
mem[16'h5E44] = 8'hAD;
mem[16'h5E45] = 8'hC5;
mem[16'h5E46] = 8'h5E;
mem[16'h5E47] = 8'hF0;
mem[16'h5E48] = 8'h19;
mem[16'h5E49] = 8'hBD;
mem[16'h5E4A] = 8'h2D;
mem[16'h5E4B] = 8'h5F;
mem[16'h5E4C] = 8'h18;
mem[16'h5E4D] = 8'h69;
mem[16'h5E4E] = 8'h28;
mem[16'h5E4F] = 8'h9D;
mem[16'h5E50] = 8'h2C;
mem[16'h5E51] = 8'h5F;
mem[16'h5E52] = 8'hA9;
mem[16'h5E53] = 8'h25;
mem[16'h5E54] = 8'h9D;
mem[16'h5E55] = 8'h1E;
mem[16'h5E56] = 8'h5F;
mem[16'h5E57] = 8'h86;
mem[16'h5E58] = 8'h70;
mem[16'h5E59] = 8'h20;
mem[16'h5E5A] = 8'hC6;
mem[16'h5E5B] = 8'h5E;
mem[16'h5E5C] = 8'hAD;
mem[16'h5E5D] = 8'hC5;
mem[16'h5E5E] = 8'h5E;
mem[16'h5E5F] = 8'h4C;
mem[16'h5E60] = 8'h1C;
mem[16'h5E61] = 8'h5E;
mem[16'h5E62] = 8'h60;
mem[16'h5E63] = 8'h02;
mem[16'h5E64] = 8'hAD;
mem[16'h5E65] = 8'hB0;
mem[16'h5E66] = 8'h4A;
mem[16'h5E67] = 8'hAA;
mem[16'h5E68] = 8'hCA;
mem[16'h5E69] = 8'hA9;
mem[16'h5E6A] = 8'h4C;
mem[16'h5E6B] = 8'h9D;
mem[16'h5E6C] = 8'h1E;
mem[16'h5E6D] = 8'h5F;
mem[16'h5E6E] = 8'hA9;
mem[16'h5E6F] = 8'h23;
mem[16'h5E70] = 8'h9D;
mem[16'h5E71] = 8'h2C;
mem[16'h5E72] = 8'h5F;
mem[16'h5E73] = 8'h86;
mem[16'h5E74] = 8'h70;
mem[16'h5E75] = 8'h20;
mem[16'h5E76] = 8'hC6;
mem[16'h5E77] = 8'h5E;
mem[16'h5E78] = 8'hAD;
mem[16'h5E79] = 8'hB0;
mem[16'h5E7A] = 8'h4A;
mem[16'h5E7B] = 8'hAA;
mem[16'h5E7C] = 8'hCA;
mem[16'h5E7D] = 8'h38;
mem[16'h5E7E] = 8'hED;
mem[16'h5E7F] = 8'hC4;
mem[16'h5E80] = 8'h5E;
mem[16'h5E81] = 8'h8D;
mem[16'h5E82] = 8'hC5;
mem[16'h5E83] = 8'h5E;
mem[16'h5E84] = 8'hCA;
mem[16'h5E85] = 8'hA9;
mem[16'h5E86] = 8'h4C;
mem[16'h5E87] = 8'h9D;
mem[16'h5E88] = 8'h1E;
mem[16'h5E89] = 8'h5F;
mem[16'h5E8A] = 8'hBD;
mem[16'h5E8B] = 8'h2D;
mem[16'h5E8C] = 8'h5F;
mem[16'h5E8D] = 8'h18;
mem[16'h5E8E] = 8'h69;
mem[16'h5E8F] = 8'h12;
mem[16'h5E90] = 8'h9D;
mem[16'h5E91] = 8'h2C;
mem[16'h5E92] = 8'h5F;
mem[16'h5E93] = 8'h86;
mem[16'h5E94] = 8'h70;
mem[16'h5E95] = 8'h20;
mem[16'h5E96] = 8'hC6;
mem[16'h5E97] = 8'h5E;
mem[16'h5E98] = 8'hA6;
mem[16'h5E99] = 8'h70;
mem[16'h5E9A] = 8'hEC;
mem[16'h5E9B] = 8'hC5;
mem[16'h5E9C] = 8'h5E;
mem[16'h5E9D] = 8'hF0;
mem[16'h5E9E] = 8'h03;
mem[16'h5E9F] = 8'h4C;
mem[16'h5EA0] = 8'h84;
mem[16'h5EA1] = 8'h5E;
mem[16'h5EA2] = 8'hCA;
mem[16'h5EA3] = 8'hAD;
mem[16'h5EA4] = 8'hC5;
mem[16'h5EA5] = 8'h5E;
mem[16'h5EA6] = 8'hC9;
mem[16'h5EA7] = 8'h08;
mem[16'h5EA8] = 8'hF0;
mem[16'h5EA9] = 8'h19;
mem[16'h5EAA] = 8'hBD;
mem[16'h5EAB] = 8'h2D;
mem[16'h5EAC] = 8'h5F;
mem[16'h5EAD] = 8'h18;
mem[16'h5EAE] = 8'h69;
mem[16'h5EAF] = 8'h44;
mem[16'h5EB0] = 8'h9D;
mem[16'h5EB1] = 8'h2C;
mem[16'h5EB2] = 8'h5F;
mem[16'h5EB3] = 8'hA9;
mem[16'h5EB4] = 8'h4C;
mem[16'h5EB5] = 8'h9D;
mem[16'h5EB6] = 8'h1E;
mem[16'h5EB7] = 8'h5F;
mem[16'h5EB8] = 8'h86;
mem[16'h5EB9] = 8'h70;
mem[16'h5EBA] = 8'h20;
mem[16'h5EBB] = 8'hC6;
mem[16'h5EBC] = 8'h5E;
mem[16'h5EBD] = 8'hAD;
mem[16'h5EBE] = 8'hC5;
mem[16'h5EBF] = 8'h5E;
mem[16'h5EC0] = 8'h4C;
mem[16'h5EC1] = 8'h7B;
mem[16'h5EC2] = 8'h5E;
mem[16'h5EC3] = 8'h60;
mem[16'h5EC4] = 8'h03;
mem[16'h5EC5] = 8'h08;
mem[16'h5EC6] = 8'hA6;
mem[16'h5EC7] = 8'h70;
mem[16'h5EC8] = 8'hBD;
mem[16'h5EC9] = 8'h83;
mem[16'h5ECA] = 8'h5B;
mem[16'h5ECB] = 8'hF0;
mem[16'h5ECC] = 8'h0B;
mem[16'h5ECD] = 8'hC9;
mem[16'h5ECE] = 8'h09;
mem[16'h5ECF] = 8'hB0;
mem[16'h5ED0] = 8'h07;
mem[16'h5ED1] = 8'hA9;
mem[16'h5ED2] = 8'h08;
mem[16'h5ED3] = 8'hA0;
mem[16'h5ED4] = 8'h5F;
mem[16'h5ED5] = 8'h4C;
mem[16'h5ED6] = 8'hDC;
mem[16'h5ED7] = 8'h5E;
mem[16'h5ED8] = 8'hA9;
mem[16'h5ED9] = 8'hF2;
mem[16'h5EDA] = 8'hA0;
mem[16'h5EDB] = 8'h5E;
mem[16'h5EDC] = 8'h20;
mem[16'h5EDD] = 8'h2B;
mem[16'h5EDE] = 8'h8C;
mem[16'h5EDF] = 8'hBD;
mem[16'h5EE0] = 8'h1E;
mem[16'h5EE1] = 8'h5F;
mem[16'h5EE2] = 8'h85;
mem[16'h5EE3] = 8'h56;
mem[16'h5EE4] = 8'hBD;
mem[16'h5EE5] = 8'h2C;
mem[16'h5EE6] = 8'h5F;
mem[16'h5EE7] = 8'h85;
mem[16'h5EE8] = 8'h57;
mem[16'h5EE9] = 8'hA9;
mem[16'h5EEA] = 8'h16;
mem[16'h5EEB] = 8'h8D;
mem[16'h5EEC] = 8'h24;
mem[16'h5EED] = 8'h8C;
mem[16'h5EEE] = 8'h20;
mem[16'h5EEF] = 8'hA8;
mem[16'h5EF0] = 8'h8B;
mem[16'h5EF1] = 8'h60;
mem[16'h5EF2] = 8'h20;
mem[16'h5EF3] = 8'h01;
mem[16'h5EF4] = 8'h20;
mem[16'h5EF5] = 8'h50;
mem[16'h5EF6] = 8'h60;
mem[16'h5EF7] = 8'h17;
mem[16'h5EF8] = 8'h7C;
mem[16'h5EF9] = 8'h1F;
mem[16'h5EFA] = 8'h65;
mem[16'h5EFB] = 8'h7F;
mem[16'h5EFC] = 8'h65;
mem[16'h5EFD] = 8'h7F;
mem[16'h5EFE] = 8'h65;
mem[16'h5EFF] = 8'h7F;
mem[16'h5F00] = 8'h7C;
mem[16'h5F01] = 8'h1F;
mem[16'h5F02] = 8'h60;
mem[16'h5F03] = 8'h17;
mem[16'h5F04] = 8'h20;
mem[16'h5F05] = 8'h50;
mem[16'h5F06] = 8'h20;
mem[16'h5F07] = 8'h01;
mem[16'h5F08] = 8'h20;
mem[16'h5F09] = 8'h00;
mem[16'h5F0A] = 8'h20;
mem[16'h5F0B] = 8'h10;
mem[16'h5F0C] = 8'h60;
mem[16'h5F0D] = 8'h17;
mem[16'h5F0E] = 8'h7C;
mem[16'h5F0F] = 8'h1F;
mem[16'h5F10] = 8'h65;
mem[16'h5F11] = 8'h7F;
mem[16'h5F12] = 8'h65;
mem[16'h5F13] = 8'h7F;
mem[16'h5F14] = 8'h65;
mem[16'h5F15] = 8'h7F;
mem[16'h5F16] = 8'h7C;
mem[16'h5F17] = 8'h1F;
mem[16'h5F18] = 8'h60;
mem[16'h5F19] = 8'h17;
mem[16'h5F1A] = 8'h20;
mem[16'h5F1B] = 8'h10;
mem[16'h5F1C] = 8'h20;
mem[16'h5F1D] = 8'h00;
mem[16'h5F1E] = 8'h25;
mem[16'h5F1F] = 8'h25;
mem[16'h5F20] = 8'h25;
mem[16'h5F21] = 8'h25;
mem[16'h5F22] = 8'h25;
mem[16'h5F23] = 8'h25;
mem[16'h5F24] = 8'h25;
mem[16'h5F25] = 8'h25;
mem[16'h5F26] = 8'h4C;
mem[16'h5F27] = 8'h4C;
mem[16'h5F28] = 8'h4C;
mem[16'h5F29] = 8'h4C;
mem[16'h5F2A] = 8'h4C;
mem[16'h5F2B] = 8'h4C;
mem[16'h5F2C] = 8'hC3;
mem[16'h5F2D] = 8'hB1;
mem[16'h5F2E] = 8'h89;
mem[16'h5F2F] = 8'h77;
mem[16'h5F30] = 8'h4F;
mem[16'h5F31] = 8'h3D;
mem[16'h5F32] = 8'h15;
mem[16'h5F33] = 8'h03;
mem[16'h5F34] = 8'hAF;
mem[16'h5F35] = 8'h9D;
mem[16'h5F36] = 8'h8B;
mem[16'h5F37] = 8'h47;
mem[16'h5F38] = 8'h35;
mem[16'h5F39] = 8'h23;
mem[16'h5F3A] = 8'hAE;
mem[16'h5F3B] = 8'hAD;
mem[16'h5F3C] = 8'h4A;
mem[16'h5F3D] = 8'h8A;
mem[16'h5F3E] = 8'h38;
mem[16'h5F3F] = 8'hE9;
mem[16'h5F40] = 8'h01;
mem[16'h5F41] = 8'h85;
mem[16'h5F42] = 8'h6E;
mem[16'h5F43] = 8'hCA;
mem[16'h5F44] = 8'h30;
mem[16'h5F45] = 8'h24;
mem[16'h5F46] = 8'h86;
mem[16'h5F47] = 8'h70;
mem[16'h5F48] = 8'hA9;
mem[16'h5F49] = 8'h7A;
mem[16'h5F4A] = 8'h9D;
mem[16'h5F4B] = 8'hB3;
mem[16'h5F4C] = 8'h60;
mem[16'h5F4D] = 8'hE4;
mem[16'h5F4E] = 8'h6E;
mem[16'h5F4F] = 8'h90;
mem[16'h5F50] = 8'h08;
mem[16'h5F51] = 8'hA9;
mem[16'h5F52] = 8'h0A;
mem[16'h5F53] = 8'h9D;
mem[16'h5F54] = 8'hAF;
mem[16'h5F55] = 8'h60;
mem[16'h5F56] = 8'h4C;
mem[16'h5F57] = 8'h62;
mem[16'h5F58] = 8'h5F;
mem[16'h5F59] = 8'hBD;
mem[16'h5F5A] = 8'hB0;
mem[16'h5F5B] = 8'h60;
mem[16'h5F5C] = 8'h18;
mem[16'h5F5D] = 8'h69;
mem[16'h5F5E] = 8'h49;
mem[16'h5F5F] = 8'h9D;
mem[16'h5F60] = 8'hAF;
mem[16'h5F61] = 8'h60;
mem[16'h5F62] = 8'h20;
mem[16'h5F63] = 8'h4D;
mem[16'h5F64] = 8'h60;
mem[16'h5F65] = 8'hA6;
mem[16'h5F66] = 8'h70;
mem[16'h5F67] = 8'h4C;
mem[16'h5F68] = 8'h43;
mem[16'h5F69] = 8'h5F;
mem[16'h5F6A] = 8'h60;
mem[16'h5F6B] = 8'hAE;
mem[16'h5F6C] = 8'hAA;
mem[16'h5F6D] = 8'h4A;
mem[16'h5F6E] = 8'h8A;
mem[16'h5F6F] = 8'h38;
mem[16'h5F70] = 8'hE9;
mem[16'h5F71] = 8'h01;
mem[16'h5F72] = 8'h85;
mem[16'h5F73] = 8'h6E;
mem[16'h5F74] = 8'hCA;
mem[16'h5F75] = 8'h30;
mem[16'h5F76] = 8'h24;
mem[16'h5F77] = 8'h86;
mem[16'h5F78] = 8'h70;
mem[16'h5F79] = 8'hA9;
mem[16'h5F7A] = 8'h95;
mem[16'h5F7B] = 8'h9D;
mem[16'h5F7C] = 8'hAB;
mem[16'h5F7D] = 8'h60;
mem[16'h5F7E] = 8'hE4;
mem[16'h5F7F] = 8'h6E;
mem[16'h5F80] = 8'h90;
mem[16'h5F81] = 8'h08;
mem[16'h5F82] = 8'hA9;
mem[16'h5F83] = 8'h0A;
mem[16'h5F84] = 8'h9D;
mem[16'h5F85] = 8'hA7;
mem[16'h5F86] = 8'h60;
mem[16'h5F87] = 8'h4C;
mem[16'h5F88] = 8'h93;
mem[16'h5F89] = 8'h5F;
mem[16'h5F8A] = 8'hBD;
mem[16'h5F8B] = 8'hA8;
mem[16'h5F8C] = 8'h60;
mem[16'h5F8D] = 8'h18;
mem[16'h5F8E] = 8'h69;
mem[16'h5F8F] = 8'h49;
mem[16'h5F90] = 8'h9D;
mem[16'h5F91] = 8'hA7;
mem[16'h5F92] = 8'h60;
mem[16'h5F93] = 8'h20;
mem[16'h5F94] = 8'h69;
mem[16'h5F95] = 8'h60;
mem[16'h5F96] = 8'hA6;
mem[16'h5F97] = 8'h70;
mem[16'h5F98] = 8'h4C;
mem[16'h5F99] = 8'h74;
mem[16'h5F9A] = 8'h5F;
mem[16'h5F9B] = 8'h60;
mem[16'h5F9C] = 8'hAE;
mem[16'h5F9D] = 8'hAC;
mem[16'h5F9E] = 8'h4A;
mem[16'h5F9F] = 8'hCA;
mem[16'h5FA0] = 8'h30;
mem[16'h5FA1] = 8'h27;
mem[16'h5FA2] = 8'h86;
mem[16'h5FA3] = 8'h70;
mem[16'h5FA4] = 8'hA9;
mem[16'h5FA5] = 8'hA3;
mem[16'h5FA6] = 8'h9D;
mem[16'h5FA7] = 8'h2E;
mem[16'h5FA8] = 8'h61;
mem[16'h5FA9] = 8'hE8;
mem[16'h5FAA] = 8'hEC;
mem[16'h5FAB] = 8'hAC;
mem[16'h5FAC] = 8'h4A;
mem[16'h5FAD] = 8'hCA;
mem[16'h5FAE] = 8'h90;
mem[16'h5FAF] = 8'h08;
mem[16'h5FB0] = 8'hA9;
mem[16'h5FB1] = 8'h1C;
mem[16'h5FB2] = 8'h9D;
mem[16'h5FB3] = 8'h2A;
mem[16'h5FB4] = 8'h61;
mem[16'h5FB5] = 8'h4C;
mem[16'h5FB6] = 8'hC1;
mem[16'h5FB7] = 8'h5F;
mem[16'h5FB8] = 8'hBD;
mem[16'h5FB9] = 8'h2B;
mem[16'h5FBA] = 8'h61;
mem[16'h5FBB] = 8'h18;
mem[16'h5FBC] = 8'h69;
mem[16'h5FBD] = 8'h62;
mem[16'h5FBE] = 8'h9D;
mem[16'h5FBF] = 8'h2A;
mem[16'h5FC0] = 8'h61;
mem[16'h5FC1] = 8'h20;
mem[16'h5FC2] = 8'hF3;
mem[16'h5FC3] = 8'h60;
mem[16'h5FC4] = 8'hA6;
mem[16'h5FC5] = 8'h70;
mem[16'h5FC6] = 8'h4C;
mem[16'h5FC7] = 8'h9F;
mem[16'h5FC8] = 8'h5F;
mem[16'h5FC9] = 8'h60;
mem[16'h5FCA] = 8'hAD;
mem[16'h5FCB] = 8'h3E;
mem[16'h5FCC] = 8'h6A;
mem[16'h5FCD] = 8'h20;
mem[16'h5FCE] = 8'h03;
mem[16'h5FCF] = 8'h9C;
mem[16'h5FD0] = 8'hC9;
mem[16'h5FD1] = 8'hA0;
mem[16'h5FD2] = 8'hF0;
mem[16'h5FD3] = 8'h0B;
mem[16'h5FD4] = 8'hC9;
mem[16'h5FD5] = 8'hC4;
mem[16'h5FD6] = 8'hD0;
mem[16'h5FD7] = 8'h08;
mem[16'h5FD8] = 8'hA9;
mem[16'h5FD9] = 8'h00;
mem[16'h5FDA] = 8'h85;
mem[16'h5FDB] = 8'h85;
mem[16'h5FDC] = 8'h20;
mem[16'h5FDD] = 8'h23;
mem[16'h5FDE] = 8'h70;
mem[16'h5FDF] = 8'h60;
mem[16'h5FE0] = 8'hC9;
mem[16'h5FE1] = 8'hCA;
mem[16'h5FE2] = 8'hD0;
mem[16'h5FE3] = 8'hE9;
mem[16'h5FE4] = 8'h85;
mem[16'h5FE5] = 8'h85;
mem[16'h5FE6] = 8'hAD;
mem[16'h5FE7] = 8'hCF;
mem[16'h5FE8] = 8'h5F;
mem[16'h5FE9] = 8'h49;
mem[16'h5FEA] = 8'h2F;
mem[16'h5FEB] = 8'h18;
mem[16'h5FEC] = 8'hC9;
mem[16'h5FED] = 8'hB1;
mem[16'h5FEE] = 8'hD0;
mem[16'h5FEF] = 8'h09;
mem[16'h5FF0] = 8'hA9;
mem[16'h5FF1] = 8'h76;
mem[16'h5FF2] = 8'h85;
mem[16'h5FF3] = 8'h89;
mem[16'h5FF4] = 8'hA9;
mem[16'h5FF5] = 8'h8A;
mem[16'h5FF6] = 8'h85;
mem[16'h5FF7] = 8'h8A;
mem[16'h5FF8] = 8'h60;
mem[16'h5FF9] = 8'hC9;
mem[16'h5FFA] = 8'hB2;
mem[16'h5FFB] = 8'hD0;
mem[16'h5FFC] = 8'h09;
mem[16'h5FFD] = 8'hA9;
mem[16'h5FFE] = 8'h6C;
mem[16'h5FFF] = 8'h85;
mem[16'h6000] = 8'h89;
mem[16'h6001] = 8'hA9;
mem[16'h6002] = 8'h94;
mem[16'h6003] = 8'h85;
mem[16'h6004] = 8'h8A;
mem[16'h6005] = 8'h60;
mem[16'h6006] = 8'hC9;
mem[16'h6007] = 8'hB3;
mem[16'h6008] = 8'hD0;
mem[16'h6009] = 8'hDF;
mem[16'h600A] = 8'hA9;
mem[16'h600B] = 8'h62;
mem[16'h600C] = 8'h85;
mem[16'h600D] = 8'h89;
mem[16'h600E] = 8'hA9;
mem[16'h600F] = 8'h9E;
mem[16'h6010] = 8'h85;
mem[16'h6011] = 8'h8A;
mem[16'h6012] = 8'h60;
mem[16'h6013] = 8'hA9;
mem[16'h6014] = 8'h2F;
mem[16'h6015] = 8'hA0;
mem[16'h6016] = 8'h60;
mem[16'h6017] = 8'h20;
mem[16'h6018] = 8'h86;
mem[16'h6019] = 8'h68;
mem[16'h601A] = 8'hA6;
mem[16'h601B] = 8'h70;
mem[16'h601C] = 8'hBD;
mem[16'h601D] = 8'h4A;
mem[16'h601E] = 8'h60;
mem[16'h601F] = 8'h85;
mem[16'h6020] = 8'h56;
mem[16'h6021] = 8'hBD;
mem[16'h6022] = 8'h47;
mem[16'h6023] = 8'h60;
mem[16'h6024] = 8'h85;
mem[16'h6025] = 8'h57;
mem[16'h6026] = 8'hA9;
mem[16'h6027] = 8'h18;
mem[16'h6028] = 8'h8D;
mem[16'h6029] = 8'h7F;
mem[16'h602A] = 8'h68;
mem[16'h602B] = 8'h20;
mem[16'h602C] = 8'hE6;
mem[16'h602D] = 8'h67;
mem[16'h602E] = 8'h60;
mem[16'h602F] = 8'h00;
mem[16'h6030] = 8'h03;
mem[16'h6031] = 8'h0C;
mem[16'h6032] = 8'h1E;
mem[16'h6033] = 8'h55;
mem[16'h6034] = 8'h0A;
mem[16'h6035] = 8'h1D;
mem[16'h6036] = 8'h55;
mem[16'h6037] = 8'h0A;
mem[16'h6038] = 8'h7D;
mem[16'h6039] = 8'h55;
mem[16'h603A] = 8'h0A;
mem[16'h603B] = 8'h7D;
mem[16'h603C] = 8'h55;
mem[16'h603D] = 8'h0A;
mem[16'h603E] = 8'h1D;
mem[16'h603F] = 8'h55;
mem[16'h6040] = 8'h0A;
mem[16'h6041] = 8'h1E;
mem[16'h6042] = 8'h55;
mem[16'h6043] = 8'h0A;
mem[16'h6044] = 8'h00;
mem[16'h6045] = 8'h03;
mem[16'h6046] = 8'h0C;
mem[16'h6047] = 8'h70;
mem[16'h6048] = 8'h0E;
mem[16'h6049] = 8'h20;
mem[16'h604A] = 8'h6C;
mem[16'h604B] = 8'h6C;
mem[16'h604C] = 8'hCB;
mem[16'h604D] = 8'hA9;
mem[16'h604E] = 8'h85;
mem[16'h604F] = 8'hA0;
mem[16'h6050] = 8'h60;
mem[16'h6051] = 8'h20;
mem[16'h6052] = 8'h2B;
mem[16'h6053] = 8'h8C;
mem[16'h6054] = 8'hA6;
mem[16'h6055] = 8'h70;
mem[16'h6056] = 8'hBD;
mem[16'h6057] = 8'hB3;
mem[16'h6058] = 8'h60;
mem[16'h6059] = 8'h85;
mem[16'h605A] = 8'h56;
mem[16'h605B] = 8'hBD;
mem[16'h605C] = 8'hAF;
mem[16'h605D] = 8'h60;
mem[16'h605E] = 8'h85;
mem[16'h605F] = 8'h57;
mem[16'h6060] = 8'hA9;
mem[16'h6061] = 8'h10;
mem[16'h6062] = 8'h8D;
mem[16'h6063] = 8'h24;
mem[16'h6064] = 8'h8C;
mem[16'h6065] = 8'h20;
mem[16'h6066] = 8'hA8;
mem[16'h6067] = 8'h8B;
mem[16'h6068] = 8'h60;
mem[16'h6069] = 8'hA9;
mem[16'h606A] = 8'h95;
mem[16'h606B] = 8'hA0;
mem[16'h606C] = 8'h60;
mem[16'h606D] = 8'h20;
mem[16'h606E] = 8'h2B;
mem[16'h606F] = 8'h8C;
mem[16'h6070] = 8'hA6;
mem[16'h6071] = 8'h70;
mem[16'h6072] = 8'hBD;
mem[16'h6073] = 8'hAB;
mem[16'h6074] = 8'h60;
mem[16'h6075] = 8'h85;
mem[16'h6076] = 8'h56;
mem[16'h6077] = 8'hBD;
mem[16'h6078] = 8'hA7;
mem[16'h6079] = 8'h60;
mem[16'h607A] = 8'h85;
mem[16'h607B] = 8'h57;
mem[16'h607C] = 8'hA9;
mem[16'h607D] = 8'h12;
mem[16'h607E] = 8'h8D;
mem[16'h607F] = 8'h24;
mem[16'h6080] = 8'h8C;
mem[16'h6081] = 8'h20;
mem[16'h6082] = 8'hA8;
mem[16'h6083] = 8'h8B;
mem[16'h6084] = 8'h60;
mem[16'h6085] = 8'h8E;
mem[16'h6086] = 8'h38;
mem[16'h6087] = 8'h8E;
mem[16'h6088] = 8'h38;
mem[16'h6089] = 8'hC4;
mem[16'h608A] = 8'h12;
mem[16'h608B] = 8'hD4;
mem[16'h608C] = 8'h2A;
mem[16'h608D] = 8'hD7;
mem[16'h608E] = 8'h2A;
mem[16'h608F] = 8'hC4;
mem[16'h6090] = 8'h12;
mem[16'h6091] = 8'h8E;
mem[16'h6092] = 8'h38;
mem[16'h6093] = 8'h8E;
mem[16'h6094] = 8'h38;
mem[16'h6095] = 8'hDB;
mem[16'h6096] = 8'h01;
mem[16'h6097] = 8'hDB;
mem[16'h6098] = 8'h21;
mem[16'h6099] = 8'hD5;
mem[16'h609A] = 8'h12;
mem[16'h609B] = 8'hD5;
mem[16'h609C] = 8'h1E;
mem[16'h609D] = 8'hD5;
mem[16'h609E] = 8'h12;
mem[16'h609F] = 8'hD5;
mem[16'h60A0] = 8'h1E;
mem[16'h60A1] = 8'hD5;
mem[16'h60A2] = 8'h12;
mem[16'h60A3] = 8'hDB;
mem[16'h60A4] = 8'h21;
mem[16'h60A5] = 8'hDB;
mem[16'h60A6] = 8'h01;
mem[16'h60A7] = 8'h9C;
mem[16'h60A8] = 8'h53;
mem[16'h60A9] = 8'h0A;
mem[16'h60AA] = 8'h20;
mem[16'h60AB] = 8'h95;
mem[16'h60AC] = 8'h95;
mem[16'h60AD] = 8'h95;
mem[16'h60AE] = 8'h0D;
mem[16'h60AF] = 8'h0A;
mem[16'h60B0] = 8'h3B;
mem[16'h60B1] = 8'h0D;
mem[16'h60B2] = 8'h0D;
mem[16'h60B3] = 8'h7A;
mem[16'h60B4] = 8'h4C;
mem[16'h60B5] = 8'h4F;
mem[16'h60B6] = 8'h47;
mem[16'h60B7] = 8'hA9;
mem[16'h60B8] = 8'hD3;
mem[16'h60B9] = 8'hA0;
mem[16'h60BA] = 8'h60;
mem[16'h60BB] = 8'h20;
mem[16'h60BC] = 8'h86;
mem[16'h60BD] = 8'h68;
mem[16'h60BE] = 8'hA6;
mem[16'h60BF] = 8'h70;
mem[16'h60C0] = 8'hBD;
mem[16'h60C1] = 8'hEF;
mem[16'h60C2] = 8'h60;
mem[16'h60C3] = 8'h85;
mem[16'h60C4] = 8'h56;
mem[16'h60C5] = 8'hBD;
mem[16'h60C6] = 8'hEB;
mem[16'h60C7] = 8'h60;
mem[16'h60C8] = 8'h85;
mem[16'h60C9] = 8'h57;
mem[16'h60CA] = 8'hA9;
mem[16'h60CB] = 8'h18;
mem[16'h60CC] = 8'h8D;
mem[16'h60CD] = 8'h7F;
mem[16'h60CE] = 8'h68;
mem[16'h60CF] = 8'h20;
mem[16'h60D0] = 8'hE6;
mem[16'h60D1] = 8'h67;
mem[16'h60D2] = 8'h60;
mem[16'h60D3] = 8'h78;
mem[16'h60D4] = 8'h30;
mem[16'h60D5] = 8'h01;
mem[16'h60D6] = 8'h54;
mem[16'h60D7] = 8'h2A;
mem[16'h60D8] = 8'h03;
mem[16'h60D9] = 8'h56;
mem[16'h60DA] = 8'h2A;
mem[16'h60DB] = 8'h0F;
mem[16'h60DC] = 8'h55;
mem[16'h60DD] = 8'h28;
mem[16'h60DE] = 8'h03;
mem[16'h60DF] = 8'h55;
mem[16'h60E0] = 8'h28;
mem[16'h60E1] = 8'h03;
mem[16'h60E2] = 8'h56;
mem[16'h60E3] = 8'h2A;
mem[16'h60E4] = 8'h0F;
mem[16'h60E5] = 8'h54;
mem[16'h60E6] = 8'h2A;
mem[16'h60E7] = 8'h03;
mem[16'h60E8] = 8'h78;
mem[16'h60E9] = 8'h30;
mem[16'h60EA] = 8'h01;
mem[16'h60EB] = 8'hCB;
mem[16'h60EC] = 8'h77;
mem[16'h60ED] = 8'h23;
mem[16'h60EE] = 8'h09;
mem[16'h60EF] = 8'h87;
mem[16'h60F0] = 8'h87;
mem[16'h60F1] = 8'h87;
mem[16'h60F2] = 8'h4C;
mem[16'h60F3] = 8'hA9;
mem[16'h60F4] = 8'h0F;
mem[16'h60F5] = 8'hA0;
mem[16'h60F6] = 8'h61;
mem[16'h60F7] = 8'h20;
mem[16'h60F8] = 8'h86;
mem[16'h60F9] = 8'h68;
mem[16'h60FA] = 8'hA6;
mem[16'h60FB] = 8'h70;
mem[16'h60FC] = 8'hBD;
mem[16'h60FD] = 8'h2E;
mem[16'h60FE] = 8'h61;
mem[16'h60FF] = 8'h85;
mem[16'h6100] = 8'h56;
mem[16'h6101] = 8'hBD;
mem[16'h6102] = 8'h2A;
mem[16'h6103] = 8'h61;
mem[16'h6104] = 8'h85;
mem[16'h6105] = 8'h57;
mem[16'h6106] = 8'hA9;
mem[16'h6107] = 8'h1B;
mem[16'h6108] = 8'h8D;
mem[16'h6109] = 8'h7F;
mem[16'h610A] = 8'h68;
mem[16'h610B] = 8'h20;
mem[16'h610C] = 8'hE6;
mem[16'h610D] = 8'h67;
mem[16'h610E] = 8'h60;
mem[16'h610F] = 8'h0F;
mem[16'h6110] = 8'h40;
mem[16'h6111] = 8'h07;
mem[16'h6112] = 8'h4F;
mem[16'h6113] = 8'h4A;
mem[16'h6114] = 8'h07;
mem[16'h6115] = 8'h56;
mem[16'h6116] = 8'h2A;
mem[16'h6117] = 8'h03;
mem[16'h6118] = 8'h15;
mem[16'h6119] = 8'h28;
mem[16'h611A] = 8'h1D;
mem[16'h611B] = 8'h15;
mem[16'h611C] = 8'h28;
mem[16'h611D] = 8'h01;
mem[16'h611E] = 8'h15;
mem[16'h611F] = 8'h28;
mem[16'h6120] = 8'h1D;
mem[16'h6121] = 8'h56;
mem[16'h6122] = 8'h2A;
mem[16'h6123] = 8'h03;
mem[16'h6124] = 8'h4F;
mem[16'h6125] = 8'h4A;
mem[16'h6126] = 8'h07;
mem[16'h6127] = 8'h0F;
mem[16'h6128] = 8'h40;
mem[16'h6129] = 8'h07;
mem[16'h612A] = 8'hE0;
mem[16'h612B] = 8'h7E;
mem[16'h612C] = 8'h1C;
mem[16'h612D] = 8'h44;
mem[16'h612E] = 8'hA3;
mem[16'h612F] = 8'hA3;
mem[16'h6130] = 8'hA3;
mem[16'h6131] = 8'h01;
mem[16'h6132] = 8'h20;
mem[16'h6133] = 8'h04;
mem[16'h6134] = 8'h00;
mem[16'h6135] = 8'h00;
mem[16'h6136] = 8'h20;
mem[16'h6137] = 8'h11;
mem[16'h6138] = 8'h02;
mem[16'h6139] = 8'h00;
mem[16'h613A] = 8'h60;
mem[16'h613B] = 8'h48;
mem[16'h613C] = 8'h00;
mem[16'h613D] = 8'h00;
mem[16'h613E] = 8'h0C;
mem[16'h613F] = 8'h60;
mem[16'h6140] = 8'h00;
mem[16'h6141] = 8'h00;
mem[16'h6142] = 8'h71;
mem[16'h6143] = 8'h00;
mem[16'h6144] = 8'h03;
mem[16'h6145] = 8'h00;
mem[16'h6146] = 8'h71;
mem[16'h6147] = 8'h00;
mem[16'h6148] = 8'h03;
mem[16'h6149] = 8'h00;
mem[16'h614A] = 8'h71;
mem[16'h614B] = 8'h00;
mem[16'h614C] = 8'h03;
mem[16'h614D] = 8'h00;
mem[16'h614E] = 8'h0C;
mem[16'h614F] = 8'h60;
mem[16'h6150] = 8'h00;
mem[16'h6151] = 8'h00;
mem[16'h6152] = 8'h60;
mem[16'h6153] = 8'h48;
mem[16'h6154] = 8'h00;
mem[16'h6155] = 8'h00;
mem[16'h6156] = 8'h20;
mem[16'h6157] = 8'h11;
mem[16'h6158] = 8'h02;
mem[16'h6159] = 8'h00;
mem[16'h615A] = 8'h20;
mem[16'h615B] = 8'h04;
mem[16'h615C] = 8'h00;
mem[16'h615D] = 8'h00;
mem[16'h615E] = 8'h40;
mem[16'h615F] = 8'h08;
mem[16'h6160] = 8'h00;
mem[16'h6161] = 8'h00;
mem[16'h6162] = 8'h40;
mem[16'h6163] = 8'h22;
mem[16'h6164] = 8'h04;
mem[16'h6165] = 8'h00;
mem[16'h6166] = 8'h40;
mem[16'h6167] = 8'h11;
mem[16'h6168] = 8'h01;
mem[16'h6169] = 8'h00;
mem[16'h616A] = 8'h18;
mem[16'h616B] = 8'h40;
mem[16'h616C] = 8'h01;
mem[16'h616D] = 8'h00;
mem[16'h616E] = 8'h62;
mem[16'h616F] = 8'h01;
mem[16'h6170] = 8'h06;
mem[16'h6171] = 8'h00;
mem[16'h6172] = 8'h62;
mem[16'h6173] = 8'h01;
mem[16'h6174] = 8'h06;
mem[16'h6175] = 8'h00;
mem[16'h6176] = 8'h62;
mem[16'h6177] = 8'h01;
mem[16'h6178] = 8'h06;
mem[16'h6179] = 8'h00;
mem[16'h617A] = 8'h18;
mem[16'h617B] = 8'h40;
mem[16'h617C] = 8'h01;
mem[16'h617D] = 8'h00;
mem[16'h617E] = 8'h40;
mem[16'h617F] = 8'h11;
mem[16'h6180] = 8'h01;
mem[16'h6181] = 8'h00;
mem[16'h6182] = 8'h40;
mem[16'h6183] = 8'h22;
mem[16'h6184] = 8'h04;
mem[16'h6185] = 8'h00;
mem[16'h6186] = 8'h40;
mem[16'h6187] = 8'h08;
mem[16'h6188] = 8'h00;
mem[16'h6189] = 8'h00;
mem[16'h618A] = 8'h00;
mem[16'h618B] = 8'h11;
mem[16'h618C] = 8'h00;
mem[16'h618D] = 8'h00;
mem[16'h618E] = 8'h00;
mem[16'h618F] = 8'h45;
mem[16'h6190] = 8'h08;
mem[16'h6191] = 8'h00;
mem[16'h6192] = 8'h00;
mem[16'h6193] = 8'h23;
mem[16'h6194] = 8'h02;
mem[16'h6195] = 8'h00;
mem[16'h6196] = 8'h30;
mem[16'h6197] = 8'h00;
mem[16'h6198] = 8'h03;
mem[16'h6199] = 8'h00;
mem[16'h619A] = 8'h44;
mem[16'h619B] = 8'h03;
mem[16'h619C] = 8'h0C;
mem[16'h619D] = 8'h00;
mem[16'h619E] = 8'h44;
mem[16'h619F] = 8'h03;
mem[16'h61A0] = 8'h0C;
mem[16'h61A1] = 8'h00;
mem[16'h61A2] = 8'h44;
mem[16'h61A3] = 8'h03;
mem[16'h61A4] = 8'h0C;
mem[16'h61A5] = 8'h00;
mem[16'h61A6] = 8'h30;
mem[16'h61A7] = 8'h00;
mem[16'h61A8] = 8'h03;
mem[16'h61A9] = 8'h00;
mem[16'h61AA] = 8'h00;
mem[16'h61AB] = 8'h23;
mem[16'h61AC] = 8'h02;
mem[16'h61AD] = 8'h00;
mem[16'h61AE] = 8'h00;
mem[16'h61AF] = 8'h45;
mem[16'h61B0] = 8'h08;
mem[16'h61B1] = 8'h00;
mem[16'h61B2] = 8'h00;
mem[16'h61B3] = 8'h11;
mem[16'h61B4] = 8'h00;
mem[16'h61B5] = 8'h00;
mem[16'h61B6] = 8'h00;
mem[16'h61B7] = 8'h22;
mem[16'h61B8] = 8'h00;
mem[16'h61B9] = 8'h00;
mem[16'h61BA] = 8'h00;
mem[16'h61BB] = 8'h0A;
mem[16'h61BC] = 8'h11;
mem[16'h61BD] = 8'h00;
mem[16'h61BE] = 8'h00;
mem[16'h61BF] = 8'h46;
mem[16'h61C0] = 8'h04;
mem[16'h61C1] = 8'h00;
mem[16'h61C2] = 8'h60;
mem[16'h61C3] = 8'h00;
mem[16'h61C4] = 8'h06;
mem[16'h61C5] = 8'h00;
mem[16'h61C6] = 8'h08;
mem[16'h61C7] = 8'h07;
mem[16'h61C8] = 8'h18;
mem[16'h61C9] = 8'h00;
mem[16'h61CA] = 8'h08;
mem[16'h61CB] = 8'h07;
mem[16'h61CC] = 8'h18;
mem[16'h61CD] = 8'h00;
mem[16'h61CE] = 8'h08;
mem[16'h61CF] = 8'h07;
mem[16'h61D0] = 8'h18;
mem[16'h61D1] = 8'h00;
mem[16'h61D2] = 8'h60;
mem[16'h61D3] = 8'h00;
mem[16'h61D4] = 8'h06;
mem[16'h61D5] = 8'h00;
mem[16'h61D6] = 8'h00;
mem[16'h61D7] = 8'h46;
mem[16'h61D8] = 8'h04;
mem[16'h61D9] = 8'h00;
mem[16'h61DA] = 8'h00;
mem[16'h61DB] = 8'h0A;
mem[16'h61DC] = 8'h11;
mem[16'h61DD] = 8'h00;
mem[16'h61DE] = 8'h00;
mem[16'h61DF] = 8'h22;
mem[16'h61E0] = 8'h00;
mem[16'h61E1] = 8'h00;
mem[16'h61E2] = 8'h00;
mem[16'h61E3] = 8'h44;
mem[16'h61E4] = 8'h00;
mem[16'h61E5] = 8'h00;
mem[16'h61E6] = 8'h00;
mem[16'h61E7] = 8'h14;
mem[16'h61E8] = 8'h22;
mem[16'h61E9] = 8'h00;
mem[16'h61EA] = 8'h00;
mem[16'h61EB] = 8'h0C;
mem[16'h61EC] = 8'h09;
mem[16'h61ED] = 8'h00;
mem[16'h61EE] = 8'h40;
mem[16'h61EF] = 8'h01;
mem[16'h61F0] = 8'h0C;
mem[16'h61F1] = 8'h00;
mem[16'h61F2] = 8'h10;
mem[16'h61F3] = 8'h0E;
mem[16'h61F4] = 8'h30;
mem[16'h61F5] = 8'h00;
mem[16'h61F6] = 8'h10;
mem[16'h61F7] = 8'h0E;
mem[16'h61F8] = 8'h30;
mem[16'h61F9] = 8'h00;
mem[16'h61FA] = 8'h10;
mem[16'h61FB] = 8'h0E;
mem[16'h61FC] = 8'h30;
mem[16'h61FD] = 8'h00;
mem[16'h61FE] = 8'h40;
mem[16'h61FF] = 8'h01;
mem[16'h6200] = 8'h0C;
mem[16'h6201] = 8'h00;
mem[16'h6202] = 8'h00;
mem[16'h6203] = 8'h0C;
mem[16'h6204] = 8'h09;
mem[16'h6205] = 8'h00;
mem[16'h6206] = 8'h00;
mem[16'h6207] = 8'h14;
mem[16'h6208] = 8'h22;
mem[16'h6209] = 8'h00;
mem[16'h620A] = 8'h00;
mem[16'h620B] = 8'h44;
mem[16'h620C] = 8'h00;
mem[16'h620D] = 8'h00;
mem[16'h620E] = 8'h00;
mem[16'h620F] = 8'h08;
mem[16'h6210] = 8'h01;
mem[16'h6211] = 8'h00;
mem[16'h6212] = 8'h00;
mem[16'h6213] = 8'h28;
mem[16'h6214] = 8'h44;
mem[16'h6215] = 8'h00;
mem[16'h6216] = 8'h00;
mem[16'h6217] = 8'h18;
mem[16'h6218] = 8'h12;
mem[16'h6219] = 8'h00;
mem[16'h621A] = 8'h00;
mem[16'h621B] = 8'h03;
mem[16'h621C] = 8'h18;
mem[16'h621D] = 8'h00;
mem[16'h621E] = 8'h20;
mem[16'h621F] = 8'h1C;
mem[16'h6220] = 8'h60;
mem[16'h6221] = 8'h00;
mem[16'h6222] = 8'h20;
mem[16'h6223] = 8'h1C;
mem[16'h6224] = 8'h60;
mem[16'h6225] = 8'h00;
mem[16'h6226] = 8'h20;
mem[16'h6227] = 8'h1C;
mem[16'h6228] = 8'h60;
mem[16'h6229] = 8'h00;
mem[16'h622A] = 8'h00;
mem[16'h622B] = 8'h03;
mem[16'h622C] = 8'h18;
mem[16'h622D] = 8'h00;
mem[16'h622E] = 8'h00;
mem[16'h622F] = 8'h18;
mem[16'h6230] = 8'h12;
mem[16'h6231] = 8'h00;
mem[16'h6232] = 8'h00;
mem[16'h6233] = 8'h28;
mem[16'h6234] = 8'h44;
mem[16'h6235] = 8'h00;
mem[16'h6236] = 8'h00;
mem[16'h6237] = 8'h08;
mem[16'h6238] = 8'h01;
mem[16'h6239] = 8'h00;
mem[16'h623A] = 8'h00;
mem[16'h623B] = 8'h10;
mem[16'h623C] = 8'h02;
mem[16'h623D] = 8'h00;
mem[16'h623E] = 8'h00;
mem[16'h623F] = 8'h50;
mem[16'h6240] = 8'h08;
mem[16'h6241] = 8'h01;
mem[16'h6242] = 8'h00;
mem[16'h6243] = 8'h30;
mem[16'h6244] = 8'h24;
mem[16'h6245] = 8'h00;
mem[16'h6246] = 8'h00;
mem[16'h6247] = 8'h06;
mem[16'h6248] = 8'h30;
mem[16'h6249] = 8'h00;
mem[16'h624A] = 8'h40;
mem[16'h624B] = 8'h38;
mem[16'h624C] = 8'h40;
mem[16'h624D] = 8'h01;
mem[16'h624E] = 8'h40;
mem[16'h624F] = 8'h38;
mem[16'h6250] = 8'h40;
mem[16'h6251] = 8'h01;
mem[16'h6252] = 8'h40;
mem[16'h6253] = 8'h38;
mem[16'h6254] = 8'h40;
mem[16'h6255] = 8'h01;
mem[16'h6256] = 8'h00;
mem[16'h6257] = 8'h06;
mem[16'h6258] = 8'h30;
mem[16'h6259] = 8'h00;
mem[16'h625A] = 8'h00;
mem[16'h625B] = 8'h30;
mem[16'h625C] = 8'h24;
mem[16'h625D] = 8'h00;
mem[16'h625E] = 8'h00;
mem[16'h625F] = 8'h50;
mem[16'h6260] = 8'h08;
mem[16'h6261] = 8'h01;
mem[16'h6262] = 8'h00;
mem[16'h6263] = 8'h10;
mem[16'h6264] = 8'h02;
mem[16'h6265] = 8'h00;
mem[16'h6266] = 8'h33;
mem[16'h6267] = 8'h45;
mem[16'h6268] = 8'h57;
mem[16'h6269] = 8'h69;
mem[16'h626A] = 8'h7B;
mem[16'h626B] = 8'h8D;
mem[16'h626C] = 8'h9F;
mem[16'h626D] = 8'h80;
mem[16'h626E] = 8'h80;
mem[16'h626F] = 8'h80;
mem[16'h6270] = 8'h80;
mem[16'h6271] = 8'h80;
mem[16'h6272] = 8'h80;
mem[16'h6273] = 8'h80;
mem[16'h6274] = 8'hB1;
mem[16'h6275] = 8'hCC;
mem[16'h6276] = 8'hE7;
mem[16'h6277] = 8'h02;
mem[16'h6278] = 8'h1D;
mem[16'h6279] = 8'h38;
mem[16'h627A] = 8'h53;
mem[16'h627B] = 8'h80;
mem[16'h627C] = 8'h80;
mem[16'h627D] = 8'h80;
mem[16'h627E] = 8'h81;
mem[16'h627F] = 8'h81;
mem[16'h6280] = 8'h81;
mem[16'h6281] = 8'h81;
mem[16'h6282] = 8'hA9;
mem[16'h6283] = 8'h00;
mem[16'h6284] = 8'h85;
mem[16'h6285] = 8'h70;
mem[16'h6286] = 8'hBD;
mem[16'h6287] = 8'hC8;
mem[16'h6288] = 8'h77;
mem[16'h6289] = 8'hC9;
mem[16'h628A] = 8'h33;
mem[16'h628B] = 8'hD0;
mem[16'h628C] = 8'h15;
mem[16'h628D] = 8'h8D;
mem[16'h628E] = 8'hBE;
mem[16'h628F] = 8'h62;
mem[16'h6290] = 8'hAD;
mem[16'h6291] = 8'h10;
mem[16'h6292] = 8'h51;
mem[16'h6293] = 8'h38;
mem[16'h6294] = 8'hE9;
mem[16'h6295] = 8'h15;
mem[16'h6296] = 8'h8D;
mem[16'h6297] = 8'hBC;
mem[16'h6298] = 8'h62;
mem[16'h6299] = 8'hA9;
mem[16'h629A] = 8'h01;
mem[16'h629B] = 8'h8D;
mem[16'h629C] = 8'hC2;
mem[16'h629D] = 8'h62;
mem[16'h629E] = 8'h20;
mem[16'h629F] = 8'hC4;
mem[16'h62A0] = 8'h62;
mem[16'h62A1] = 8'h60;
mem[16'h62A2] = 8'hA9;
mem[16'h62A3] = 8'hEA;
mem[16'h62A4] = 8'h8D;
mem[16'h62A5] = 8'hD8;
mem[16'h62A6] = 8'h77;
mem[16'h62A7] = 8'h8D;
mem[16'h62A8] = 8'hBC;
mem[16'h62A9] = 8'h62;
mem[16'h62AA] = 8'hA9;
mem[16'h62AB] = 8'h5E;
mem[16'h62AC] = 8'h8D;
mem[16'h62AD] = 8'hBE;
mem[16'h62AE] = 8'h62;
mem[16'h62AF] = 8'hA9;
mem[16'h62B0] = 8'h01;
mem[16'h62B1] = 8'h8D;
mem[16'h62B2] = 8'hC2;
mem[16'h62B3] = 8'h62;
mem[16'h62B4] = 8'h20;
mem[16'h62B5] = 8'hC4;
mem[16'h62B6] = 8'h62;
mem[16'h62B7] = 8'h60;
mem[16'h62B8] = 8'h20;
mem[16'h62B9] = 8'h20;
mem[16'h62BA] = 8'h20;
mem[16'h62BB] = 8'h20;
mem[16'h62BC] = 8'hE5;
mem[16'h62BD] = 8'h20;
mem[16'h62BE] = 8'h30;
mem[16'h62BF] = 8'h2C;
mem[16'h62C0] = 8'h00;
mem[16'h62C1] = 8'h00;
mem[16'h62C2] = 8'h00;
mem[16'h62C3] = 8'h00;
mem[16'h62C4] = 8'hA9;
mem[16'h62C5] = 8'hE0;
mem[16'h62C6] = 8'hA0;
mem[16'h62C7] = 8'h62;
mem[16'h62C8] = 8'h20;
mem[16'h62C9] = 8'h86;
mem[16'h62CA] = 8'h68;
mem[16'h62CB] = 8'hA9;
mem[16'h62CC] = 8'h18;
mem[16'h62CD] = 8'h8D;
mem[16'h62CE] = 8'h7F;
mem[16'h62CF] = 8'h68;
mem[16'h62D0] = 8'hA6;
mem[16'h62D1] = 8'h70;
mem[16'h62D2] = 8'hBD;
mem[16'h62D3] = 8'hBC;
mem[16'h62D4] = 8'h62;
mem[16'h62D5] = 8'h85;
mem[16'h62D6] = 8'h57;
mem[16'h62D7] = 8'hBD;
mem[16'h62D8] = 8'hBE;
mem[16'h62D9] = 8'h62;
mem[16'h62DA] = 8'h85;
mem[16'h62DB] = 8'h56;
mem[16'h62DC] = 8'h20;
mem[16'h62DD] = 8'hE6;
mem[16'h62DE] = 8'h67;
mem[16'h62DF] = 8'h60;
mem[16'h62E0] = 8'h39;
mem[16'h62E1] = 8'h00;
mem[16'h62E2] = 8'h00;
mem[16'h62E3] = 8'h6E;
mem[16'h62E4] = 8'h00;
mem[16'h62E5] = 8'h00;
mem[16'h62E6] = 8'h70;
mem[16'h62E7] = 8'h00;
mem[16'h62E8] = 8'h00;
mem[16'h62E9] = 8'h60;
mem[16'h62EA] = 8'h00;
mem[16'h62EB] = 8'h03;
mem[16'h62EC] = 8'h40;
mem[16'h62ED] = 8'h41;
mem[16'h62EE] = 8'h07;
mem[16'h62EF] = 8'h00;
mem[16'h62F0] = 8'h63;
mem[16'h62F1] = 8'h0C;
mem[16'h62F2] = 8'h00;
mem[16'h62F3] = 8'h3E;
mem[16'h62F4] = 8'h18;
mem[16'h62F5] = 8'h00;
mem[16'h62F6] = 8'h1C;
mem[16'h62F7] = 8'h10;
mem[16'h62F8] = 8'hA9;
mem[16'h62F9] = 8'h14;
mem[16'h62FA] = 8'hA0;
mem[16'h62FB] = 8'h63;
mem[16'h62FC] = 8'h20;
mem[16'h62FD] = 8'h86;
mem[16'h62FE] = 8'h68;
mem[16'h62FF] = 8'hA9;
mem[16'h6300] = 8'h18;
mem[16'h6301] = 8'h8D;
mem[16'h6302] = 8'h7F;
mem[16'h6303] = 8'h68;
mem[16'h6304] = 8'hA6;
mem[16'h6305] = 8'h70;
mem[16'h6306] = 8'hBD;
mem[16'h6307] = 8'hB8;
mem[16'h6308] = 8'h62;
mem[16'h6309] = 8'h85;
mem[16'h630A] = 8'h57;
mem[16'h630B] = 8'hBD;
mem[16'h630C] = 8'hBA;
mem[16'h630D] = 8'h62;
mem[16'h630E] = 8'h85;
mem[16'h630F] = 8'h56;
mem[16'h6310] = 8'h20;
mem[16'h6311] = 8'hE6;
mem[16'h6312] = 8'h67;
mem[16'h6313] = 8'h60;
mem[16'h6314] = 8'h00;
mem[16'h6315] = 8'h40;
mem[16'h6316] = 8'h13;
mem[16'h6317] = 8'h00;
mem[16'h6318] = 8'h60;
mem[16'h6319] = 8'h0E;
mem[16'h631A] = 8'h00;
mem[16'h631B] = 8'h60;
mem[16'h631C] = 8'h01;
mem[16'h631D] = 8'h18;
mem[16'h631E] = 8'h60;
mem[16'h631F] = 8'h00;
mem[16'h6320] = 8'h3C;
mem[16'h6321] = 8'h30;
mem[16'h6322] = 8'h00;
mem[16'h6323] = 8'h66;
mem[16'h6324] = 8'h18;
mem[16'h6325] = 8'h00;
mem[16'h6326] = 8'h43;
mem[16'h6327] = 8'h0F;
mem[16'h6328] = 8'h00;
mem[16'h6329] = 8'h01;
mem[16'h632A] = 8'h07;
mem[16'h632B] = 8'h00;
mem[16'h632C] = 8'h42;
mem[16'h632D] = 8'h47;
mem[16'h632E] = 8'h4E;
mem[16'h632F] = 8'h31;
mem[16'h6330] = 8'h0D;
mem[16'h6331] = 8'h0A;
mem[16'h6332] = 8'hCD;
mem[16'h6333] = 8'h02;
mem[16'h6334] = 8'h23;
mem[16'h6335] = 8'h4C;
mem[16'h6336] = 8'h4F;
mem[16'h6337] = 8'h47;
mem[16'h6338] = 8'h53;
mem[16'h6339] = 8'h54;
mem[16'h633A] = 8'h52;
mem[16'h633B] = 8'h0D;
mem[16'h633C] = 8'h0A;
mem[16'h633D] = 8'hCF;
mem[16'h633E] = 8'h02;
mem[16'h633F] = 8'h2F;
mem[16'h6340] = 8'h4C;
mem[16'h6341] = 8'h4F;
mem[16'h6342] = 8'h47;
mem[16'h6343] = 8'h53;
mem[16'h6344] = 8'h54;
mem[16'h6345] = 8'h52;
mem[16'h6346] = 8'h0D;
mem[16'h6347] = 8'h09;
mem[16'h6348] = 8'hCB;
mem[16'h6349] = 8'h01;
mem[16'h634A] = 8'h4E;
mem[16'h634B] = 8'h53;
mem[16'h634C] = 8'h54;
mem[16'h634D] = 8'h4F;
mem[16'h634E] = 8'h52;
mem[16'h634F] = 8'h45;
mem[16'h6350] = 8'h0D;
mem[16'h6351] = 8'h05;
mem[16'h6352] = 8'hCD;
mem[16'h6353] = 8'h02;
mem[16'h6354] = 8'h23;
mem[16'h6355] = 8'h39;
mem[16'h6356] = 8'h0D;
mem[16'h6357] = 8'h09;
mem[16'h6358] = 8'hD0;
mem[16'h6359] = 8'h01;
mem[16'h635A] = 8'h4E;
mem[16'h635B] = 8'h50;
mem[16'h635C] = 8'h4C;
mem[16'h635D] = 8'h45;
mem[16'h635E] = 8'h2B;
mem[16'h635F] = 8'h31;
mem[16'h6360] = 8'h0D;
mem[16'h6361] = 8'h08;
mem[16'h6362] = 8'hD0;
mem[16'h6363] = 8'h06;
mem[16'h6364] = 8'h42;
mem[16'h6365] = 8'h47;
mem[16'h6366] = 8'h4E;
mem[16'h6367] = 8'h2C;
mem[16'h6368] = 8'h58;
mem[16'h6369] = 8'h0D;
mem[16'h636A] = 8'h08;
mem[16'h636B] = 8'hCB;
mem[16'h636C] = 8'h01;
mem[16'h636D] = 8'h4E;
mem[16'h636E] = 8'h50;
mem[16'h636F] = 8'h4C;
mem[16'h6370] = 8'h4F;
mem[16'h6371] = 8'h54;
mem[16'h6372] = 8'h0D;
mem[16'h6373] = 8'h0F;
mem[16'h6374] = 8'h4C;
mem[16'h6375] = 8'h47;
mem[16'h6376] = 8'h42;
mem[16'h6377] = 8'h47;
mem[16'h6378] = 8'h4E;
mem[16'h6379] = 8'h31;
mem[16'h637A] = 8'h20;
mem[16'h637B] = 8'h20;
mem[16'h637C] = 8'hCE;
mem[16'h637D] = 8'h01;
mem[16'h637E] = 8'h58;
mem[16'h637F] = 8'h49;
mem[16'h6380] = 8'h4E;
mem[16'h6381] = 8'h44;
mem[16'h6382] = 8'h0D;
mem[16'h6383] = 8'h09;
mem[16'h6384] = 8'hCD;
mem[16'h6385] = 8'h06;
mem[16'h6386] = 8'h59;
mem[16'h6387] = 8'h4C;
mem[16'h6388] = 8'h4F;
mem[16'h6389] = 8'h47;
mem[16'h638A] = 8'h2C;
mem[16'h638B] = 8'h58;
mem[16'h638C] = 8'h0D;
mem[16'h638D] = 8'h08;
mem[16'h638E] = 8'hD0;
mem[16'h638F] = 8'h01;
mem[16'h6390] = 8'h59;
mem[16'h6391] = 8'h41;
mem[16'h6392] = 8'h58;
mem[16'h6393] = 8'h49;
mem[16'h6394] = 8'h53;
mem[16'h6395] = 8'h0D;
mem[16'h6396] = 8'h09;
mem[16'h6397] = 8'hCF;
mem[16'h6398] = 8'h06;
mem[16'h6399] = 8'h58;
mem[16'h639A] = 8'h4C;
mem[16'h639B] = 8'h4F;
mem[16'h639C] = 8'h47;
mem[16'h639D] = 8'h2C;
mem[16'h639E] = 8'h58;
mem[16'h639F] = 8'h0D;
mem[16'h63A0] = 8'h08;
mem[16'h63A1] = 8'hD2;
mem[16'h63A2] = 8'h01;
mem[16'h63A3] = 8'h58;
mem[16'h63A4] = 8'h41;
mem[16'h63A5] = 8'h58;
mem[16'h63A6] = 8'h49;
mem[16'h63A7] = 8'h53;
mem[16'h63A8] = 8'h0D;
mem[16'h63A9] = 8'h0B;
mem[16'h63AA] = 8'hCD;
mem[16'h63AB] = 8'h07;
mem[16'h63AC] = 8'h58;
mem[16'h63AD] = 8'h43;
mem[16'h63AE] = 8'h4F;
mem[16'h63AF] = 8'h4F;
mem[16'h63B0] = 8'h52;
mem[16'h63B1] = 8'h44;
mem[16'h63B2] = 8'h2C;
mem[16'h63B3] = 8'h59;
mem[16'h63B4] = 8'h0D;
mem[16'h63B5] = 8'h03;
mem[16'h63B6] = 8'hAC;
mem[16'h63B7] = 8'h00;
mem[16'h63B8] = 8'h0D;
mem[16'h63B9] = 8'h0B;
mem[16'h63BA] = 8'hCD;
mem[16'h63BB] = 8'h06;
mem[16'h63BC] = 8'h42;
mem[16'h63BD] = 8'h49;
mem[16'h63BE] = 8'h54;
mem[16'h63BF] = 8'h43;
mem[16'h63C0] = 8'h4E;
mem[16'h63C1] = 8'h56;
mem[16'h63C2] = 8'h2C;
mem[16'h63C3] = 8'h58;
mem[16'h63C4] = 8'h0D;
mem[16'h63C5] = 8'h03;
mem[16'h63C6] = 8'hAC;
mem[16'h63C7] = 8'h00;
mem[16'h63C8] = 8'h0D;
mem[16'h63C9] = 8'h0A;
mem[16'h63CA] = 8'hCD;
mem[16'h63CB] = 8'h06;
mem[16'h63CC] = 8'h53;
mem[16'h63CD] = 8'h43;
mem[16'h63CE] = 8'h32;
mem[16'h63CF] = 8'h4C;
mem[16'h63D0] = 8'h4F;
mem[16'h63D1] = 8'h2C;
mem[16'h63D2] = 8'h58;
mem[16'h63D3] = 8'h0D;
mem[16'h63D4] = 8'h0A;
mem[16'h63D5] = 8'hCF;
mem[16'h63D6] = 8'h06;
mem[16'h63D7] = 8'h53;
mem[16'h63D8] = 8'h43;
mem[16'h63D9] = 8'h32;
mem[16'h63DA] = 8'h48;
mem[16'h63DB] = 8'h49;
mem[16'h63DC] = 8'h2C;
mem[16'h63DD] = 8'h58;
mem[16'h63DE] = 8'h0D;
mem[16'h63DF] = 8'h09;
mem[16'h63E0] = 8'hCB;
mem[16'h63E1] = 8'h01;
mem[16'h63E2] = 8'h45;
mem[16'h63E3] = 8'h53;
mem[16'h63E4] = 8'h54;
mem[16'h63E5] = 8'h4F;
mem[16'h63E6] = 8'h52;
mem[16'h63E7] = 8'h45;
mem[16'h63E8] = 8'h0D;
mem[16'h63E9] = 8'h06;
mem[16'h63EA] = 8'hCD;
mem[16'h63EB] = 8'h02;
mem[16'h63EC] = 8'h23;
mem[16'h63ED] = 8'h31;
mem[16'h63EE] = 8'h38;
mem[16'h63EF] = 8'h0D;
mem[16'h63F0] = 8'h09;
mem[16'h63F1] = 8'hD0;
mem[16'h63F2] = 8'h01;
mem[16'h63F3] = 8'h45;
mem[16'h63F4] = 8'h50;
mem[16'h63F5] = 8'h4C;
mem[16'h63F6] = 8'h45;
mem[16'h63F7] = 8'h2B;
mem[16'h63F8] = 8'h31;
mem[16'h63F9] = 8'h0D;
mem[16'h63FA] = 8'h08;
mem[16'h63FB] = 8'hCB;
mem[16'h63FC] = 8'h01;
mem[16'h63FD] = 8'h45;
mem[16'h63FE] = 8'h50;
mem[16'h63FF] = 8'h4C;
mem[16'h6400] = 8'h4F;
mem[16'h6401] = 8'h54;
mem[16'h6402] = 8'h0D;
mem[16'h6403] = 8'h03;
mem[16'h6404] = 8'hA5;
mem[16'h6405] = 8'h00;
mem[16'h6406] = 8'h0D;
mem[16'h6407] = 8'h10;
mem[16'h6408] = 8'h4C;
mem[16'h6409] = 8'h47;
mem[16'h640A] = 8'h42;
mem[16'h640B] = 8'h47;
mem[16'h640C] = 8'h4E;
mem[16'h640D] = 8'h33;
mem[16'h640E] = 8'h20;
mem[16'h640F] = 8'h20;
mem[16'h6410] = 8'hCD;
mem[16'h6411] = 8'h06;
mem[16'h6412] = 8'h42;
mem[16'h6413] = 8'h47;
mem[16'h6414] = 8'h4E;
mem[16'h6415] = 8'h2C;
mem[16'h6416] = 8'h58;
mem[16'h6417] = 8'h0D;
mem[16'h6418] = 8'h09;
mem[16'h6419] = 8'h87;
mem[16'h641A] = 8'h01;
mem[16'h641B] = 8'h4C;
mem[16'h641C] = 8'h47;
mem[16'h641D] = 8'h42;
mem[16'h641E] = 8'h47;
mem[16'h641F] = 8'h4E;
mem[16'h6420] = 8'h34;
mem[16'h6421] = 8'h0D;
mem[16'h6422] = 8'h0A;
mem[16'h6423] = 8'hCD;
mem[16'h6424] = 8'h02;
mem[16'h6425] = 8'h23;
mem[16'h6426] = 8'h4C;
mem[16'h6427] = 8'h4F;
mem[16'h6428] = 8'h47;
mem[16'h6429] = 8'h53;
mem[16'h642A] = 8'h54;
mem[16'h642B] = 8'h52;
mem[16'h642C] = 8'h0D;
mem[16'h642D] = 8'h0A;
mem[16'h642E] = 8'hCF;
mem[16'h642F] = 8'h02;
mem[16'h6430] = 8'h2F;
mem[16'h6431] = 8'h4C;
mem[16'h6432] = 8'h4F;
mem[16'h6433] = 8'h47;
mem[16'h6434] = 8'h53;
mem[16'h6435] = 8'h54;
mem[16'h6436] = 8'h52;
mem[16'h6437] = 8'h0D;
mem[16'h6438] = 8'h09;
mem[16'h6439] = 8'hCB;
mem[16'h643A] = 8'h01;
mem[16'h643B] = 8'h4E;
mem[16'h643C] = 8'h53;
mem[16'h643D] = 8'h54;
mem[16'h643E] = 8'h4F;
mem[16'h643F] = 8'h52;
mem[16'h6440] = 8'h45;
mem[16'h6441] = 8'h0D;
mem[16'h6442] = 8'h05;
mem[16'h6443] = 8'hCD;
mem[16'h6444] = 8'h02;
mem[16'h6445] = 8'h23;
mem[16'h6446] = 8'h39;
mem[16'h6447] = 8'h0D;
mem[16'h6448] = 8'h09;
mem[16'h6449] = 8'hD0;
mem[16'h644A] = 8'h01;
mem[16'h644B] = 8'h4E;
mem[16'h644C] = 8'h50;
mem[16'h644D] = 8'h4C;
mem[16'h644E] = 8'h45;
mem[16'h644F] = 8'h2B;
mem[16'h6450] = 8'h31;
mem[16'h6451] = 8'h0D;
mem[16'h6452] = 8'h08;
mem[16'h6453] = 8'hCB;
mem[16'h6454] = 8'h01;
mem[16'h6455] = 8'h4E;
mem[16'h6456] = 8'h50;
mem[16'h6457] = 8'h4C;
mem[16'h6458] = 8'h4F;
mem[16'h6459] = 8'h54;
mem[16'h645A] = 8'h0D;
mem[16'h645B] = 8'h07;
mem[16'h645C] = 8'hCE;
mem[16'h645D] = 8'h01;
mem[16'h645E] = 8'h58;
mem[16'h645F] = 8'h49;
mem[16'h6460] = 8'h4E;
mem[16'h6461] = 8'h44;
mem[16'h6462] = 8'h0D;
mem[16'h6463] = 8'h05;
mem[16'h6464] = 8'hCD;
mem[16'h6465] = 8'h02;
mem[16'h6466] = 8'h23;
mem[16'h6467] = 8'h30;
mem[16'h6468] = 8'h0D;
mem[16'h6469] = 8'h08;
mem[16'h646A] = 8'hD0;
mem[16'h646B] = 8'h06;
mem[16'h646C] = 8'h42;
mem[16'h646D] = 8'h47;
mem[16'h646E] = 8'h4E;
mem[16'h646F] = 8'h2C;
mem[16'h6470] = 8'h58;
mem[16'h6471] = 8'h0D;
mem[16'h6472] = 8'h0B;
mem[16'h6473] = 8'h4C;
mem[16'h6474] = 8'h47;
mem[16'h6475] = 8'h42;
mem[16'h6476] = 8'h47;
mem[16'h6477] = 8'h4E;
mem[16'h6478] = 8'h34;
mem[16'h6479] = 8'h20;
mem[16'h647A] = 8'h20;
mem[16'h647B] = 8'hA5;
mem[16'h647C] = 8'h00;
mem[16'h647D] = 8'h0D;
mem[16'h647E] = 8'h03;
mem[16'h647F] = 8'h3B;
mem[16'h6480] = 8'h20;
mem[16'h6481] = 8'h0D;
mem[16'h6482] = 8'h0F;
mem[16'h6483] = 8'h4C;
mem[16'h6484] = 8'h4F;
mem[16'h6485] = 8'h47;
mem[16'h6486] = 8'h45;
mem[16'h6487] = 8'h4E;
mem[16'h6488] = 8'h44;
mem[16'h6489] = 8'h20;
mem[16'h648A] = 8'h20;
mem[16'h648B] = 8'hCE;
mem[16'h648C] = 8'h01;
mem[16'h648D] = 8'h58;
mem[16'h648E] = 8'h49;
mem[16'h648F] = 8'h4E;
mem[16'h6490] = 8'h44;
mem[16'h6491] = 8'h0D;
mem[16'h6492] = 8'h09;
mem[16'h6493] = 8'hCD;
mem[16'h6494] = 8'h06;
mem[16'h6495] = 8'h45;
mem[16'h6496] = 8'h4E;
mem[16'h6497] = 8'h44;
mem[16'h6498] = 8'h4C;
mem[16'h6499] = 8'h2C;
mem[16'h649A] = 8'h58;
mem[16'h649B] = 8'h0D;
mem[16'h649C] = 8'h0A;
mem[16'h649D] = 8'h86;
mem[16'h649E] = 8'h01;
mem[16'h649F] = 8'h4C;
mem[16'h64A0] = 8'h4F;
mem[16'h64A1] = 8'h47;
mem[16'h64A2] = 8'h45;
mem[16'h64A3] = 8'h4E;
mem[16'h64A4] = 8'h44;
mem[16'h64A5] = 8'h31;
mem[16'h64A6] = 8'h0D;
mem[16'h64A7] = 8'h0F;
mem[16'h64A8] = 8'h4C;
mem[16'h64A9] = 8'h4F;
mem[16'h64AA] = 8'h47;
mem[16'h64AB] = 8'h45;
mem[16'h64AC] = 8'h4E;
mem[16'h64AD] = 8'h44;
mem[16'h64AE] = 8'h30;
mem[16'h64AF] = 8'h20;
mem[16'h64B0] = 8'hCE;
mem[16'h64B1] = 8'h01;
mem[16'h64B2] = 8'h58;
mem[16'h64B3] = 8'h49;
mem[16'h64B4] = 8'h4E;
mem[16'h64B5] = 8'h44;
mem[16'h64B6] = 8'h0D;
mem[16'h64B7] = 8'h09;
mem[16'h64B8] = 8'hCD;
mem[16'h64B9] = 8'h06;
mem[16'h64BA] = 8'h59;
mem[16'h64BB] = 8'h4C;
mem[16'h64BC] = 8'h4F;
mem[16'h64BD] = 8'h47;
mem[16'h64BE] = 8'h2C;
mem[16'h64BF] = 8'h58;
mem[16'h64C0] = 8'h0D;
mem[16'h64C1] = 8'h08;
mem[16'h64C2] = 8'hD0;
mem[16'h64C3] = 8'h01;
mem[16'h64C4] = 8'h59;
mem[16'h64C5] = 8'h41;
mem[16'h64C6] = 8'h58;
mem[16'h64C7] = 8'h49;
mem[16'h64C8] = 8'h53;
mem[16'h64C9] = 8'h0D;
mem[16'h64CA] = 8'h09;
mem[16'h64CB] = 8'hCD;
mem[16'h64CC] = 8'h06;
mem[16'h64CD] = 8'h58;
mem[16'h64CE] = 8'h4C;
mem[16'h64CF] = 8'h4F;
mem[16'h64D0] = 8'h47;
mem[16'h64D1] = 8'h2C;
mem[16'h64D2] = 8'h58;
mem[16'h64D3] = 8'h0D;
mem[16'h64D4] = 8'h03;
mem[16'h64D5] = 8'hA9;
mem[16'h64D6] = 8'h00;
mem[16'h64D7] = 8'h0D;
mem[16'h64D8] = 8'h0B;
mem[16'h64D9] = 8'hF0;
mem[16'h64DA] = 8'h06;
mem[16'h64DB] = 8'h4C;
mem[16'h64DC] = 8'h45;
mem[16'h64DD] = 8'h4E;
mem[16'h64DE] = 8'h4C;
mem[16'h64DF] = 8'h4F;
mem[16'h64E0] = 8'h47;
mem[16'h64E1] = 8'h2C;
mem[16'h64E2] = 8'h58;
mem[16'h64E3] = 8'h0D;
mem[16'h64E4] = 8'h0A;
mem[16'h64E5] = 8'h83;
mem[16'h64E6] = 8'h01;
mem[16'h64E7] = 8'h4C;
mem[16'h64E8] = 8'h4F;
mem[16'h64E9] = 8'h47;
mem[16'h64EA] = 8'h45;
mem[16'h64EB] = 8'h4E;
mem[16'h64EC] = 8'h44;
mem[16'h64ED] = 8'h31;
mem[16'h64EE] = 8'h0D;
mem[16'h64EF] = 8'h08;
mem[16'h64F0] = 8'hD0;
mem[16'h64F1] = 8'h01;
mem[16'h64F2] = 8'h58;
mem[16'h64F3] = 8'h41;
mem[16'h64F4] = 8'h58;
mem[16'h64F5] = 8'h49;
mem[16'h64F6] = 8'h53;
mem[16'h64F7] = 8'h0D;
mem[16'h64F8] = 8'h05;
mem[16'h64F9] = 8'hCD;
mem[16'h64FA] = 8'h02;
mem[16'h64FB] = 8'h23;
mem[16'h64FC] = 8'h39;
mem[16'h64FD] = 8'h0D;
mem[16'h64FE] = 8'h09;
mem[16'h64FF] = 8'hD0;
mem[16'h6500] = 8'hA5;
mem[16'h6501] = 8'h55;
mem[16'h6502] = 8'h29;
mem[16'h6503] = 8'h7F;
mem[16'h6504] = 8'hA8;
mem[16'h6505] = 8'hA6;
mem[16'h6506] = 8'h50;
mem[16'h6507] = 8'hAD;
mem[16'h6508] = 8'h30;
mem[16'h6509] = 8'hC0;
mem[16'h650A] = 8'hCA;
mem[16'h650B] = 8'hD0;
mem[16'h650C] = 8'h05;
mem[16'h650D] = 8'hA6;
mem[16'h650E] = 8'h50;
mem[16'h650F] = 8'hAD;
mem[16'h6510] = 8'h30;
mem[16'h6511] = 8'hC0;
mem[16'h6512] = 8'hA5;
mem[16'h6513] = 8'h55;
mem[16'h6514] = 8'hF0;
mem[16'h6515] = 8'h10;
mem[16'h6516] = 8'h88;
mem[16'h6517] = 8'hD0;
mem[16'h6518] = 8'h0D;
mem[16'h6519] = 8'hA8;
mem[16'h651A] = 8'h30;
mem[16'h651B] = 8'h05;
mem[16'h651C] = 8'hC6;
mem[16'h651D] = 8'h50;
mem[16'h651E] = 8'h98;
mem[16'h651F] = 8'hD0;
mem[16'h6520] = 8'h05;
mem[16'h6521] = 8'hE6;
mem[16'h6522] = 8'h50;
mem[16'h6523] = 8'h29;
mem[16'h6524] = 8'h7F;
mem[16'h6525] = 8'hA8;
mem[16'h6526] = 8'hC6;
mem[16'h6527] = 8'h52;
mem[16'h6528] = 8'hD0;
mem[16'h6529] = 8'hE0;
mem[16'h652A] = 8'hC6;
mem[16'h652B] = 8'h53;
mem[16'h652C] = 8'h10;
mem[16'h652D] = 8'hDC;
mem[16'h652E] = 8'h60;
mem[16'h652F] = 8'hAD;
mem[16'h6530] = 8'h54;
mem[16'h6531] = 8'hC0;
mem[16'h6532] = 8'hAD;
mem[16'h6533] = 8'h52;
mem[16'h6534] = 8'hC0;
mem[16'h6535] = 8'hAD;
mem[16'h6536] = 8'h57;
mem[16'h6537] = 8'hC0;
mem[16'h6538] = 8'hAD;
mem[16'h6539] = 8'h50;
mem[16'h653A] = 8'hC0;
mem[16'h653B] = 8'hA9;
mem[16'h653C] = 8'h00;
mem[16'h653D] = 8'h85;
mem[16'h653E] = 8'h64;
mem[16'h653F] = 8'h85;
mem[16'h6540] = 8'h65;
mem[16'h6541] = 8'h60;
mem[16'h6542] = 8'hA9;
mem[16'h6543] = 8'h00;
mem[16'h6544] = 8'h85;
mem[16'h6545] = 8'h59;
mem[16'h6546] = 8'hA9;
mem[16'h6547] = 8'h20;
mem[16'h6548] = 8'h85;
mem[16'h6549] = 8'h5A;
mem[16'h654A] = 8'hA9;
mem[16'h654B] = 8'h00;
mem[16'h654C] = 8'hA0;
mem[16'h654D] = 8'h00;
mem[16'h654E] = 8'h91;
mem[16'h654F] = 8'h59;
mem[16'h6550] = 8'hA5;
mem[16'h6551] = 8'h59;
mem[16'h6552] = 8'h18;
mem[16'h6553] = 8'h69;
mem[16'h6554] = 8'h01;
mem[16'h6555] = 8'h85;
mem[16'h6556] = 8'h59;
mem[16'h6557] = 8'hA5;
mem[16'h6558] = 8'h5A;
mem[16'h6559] = 8'h69;
mem[16'h655A] = 8'h00;
mem[16'h655B] = 8'h85;
mem[16'h655C] = 8'h5A;
mem[16'h655D] = 8'hC9;
mem[16'h655E] = 8'h40;
mem[16'h655F] = 8'hD0;
mem[16'h6560] = 8'hE9;
mem[16'h6561] = 8'h60;
mem[16'h6562] = 8'h10;
mem[16'h6563] = 8'h05;
mem[16'h6564] = 8'h49;
mem[16'h6565] = 8'hFF;
mem[16'h6566] = 8'h18;
mem[16'h6567] = 8'h69;
mem[16'h6568] = 8'h01;
mem[16'h6569] = 8'h60;
mem[16'h656A] = 8'hA2;
mem[16'h656B] = 8'h00;
mem[16'h656C] = 8'hA4;
mem[16'h656D] = 8'h56;
mem[16'h656E] = 8'hC0;
mem[16'h656F] = 8'hC0;
mem[16'h6570] = 8'hB0;
mem[16'h6571] = 8'h4A;
mem[16'h6572] = 8'hB9;
mem[16'h6573] = 8'hD5;
mem[16'h6574] = 8'h8E;
mem[16'h6575] = 8'h85;
mem[16'h6576] = 8'h59;
mem[16'h6577] = 8'hB9;
mem[16'h6578] = 8'h95;
mem[16'h6579] = 8'h8F;
mem[16'h657A] = 8'h85;
mem[16'h657B] = 8'h5A;
mem[16'h657C] = 8'hA4;
mem[16'h657D] = 8'h57;
mem[16'h657E] = 8'hB9;
mem[16'h657F] = 8'h3E;
mem[16'h6580] = 8'h8C;
mem[16'h6581] = 8'h85;
mem[16'h6582] = 8'h5C;
mem[16'h6583] = 8'hB9;
mem[16'h6584] = 8'h56;
mem[16'h6585] = 8'h8D;
mem[16'h6586] = 8'hA8;
mem[16'h6587] = 8'hBD;
mem[16'h6588] = 8'h79;
mem[16'h6589] = 8'h51;
mem[16'h658A] = 8'h29;
mem[16'h658B] = 8'h80;
mem[16'h658C] = 8'h85;
mem[16'h658D] = 8'h6D;
mem[16'h658E] = 8'hBD;
mem[16'h658F] = 8'h79;
mem[16'h6590] = 8'h51;
mem[16'h6591] = 8'h29;
mem[16'h6592] = 8'h7F;
mem[16'h6593] = 8'h85;
mem[16'h6594] = 8'h66;
mem[16'h6595] = 8'hA9;
mem[16'h6596] = 8'h00;
mem[16'h6597] = 8'h85;
mem[16'h6598] = 8'h6A;
mem[16'h6599] = 8'hA5;
mem[16'h659A] = 8'h5C;
mem[16'h659B] = 8'hC9;
mem[16'h659C] = 8'h01;
mem[16'h659D] = 8'hF0;
mem[16'h659E] = 8'h15;
mem[16'h659F] = 8'h46;
mem[16'h65A0] = 8'h66;
mem[16'h65A1] = 8'h66;
mem[16'h65A2] = 8'h6A;
mem[16'h65A3] = 8'h06;
mem[16'h65A4] = 8'h5C;
mem[16'h65A5] = 8'h24;
mem[16'h65A6] = 8'h5C;
mem[16'h65A7] = 8'h10;
mem[16'h65A8] = 8'hF6;
mem[16'h65A9] = 8'h46;
mem[16'h65AA] = 8'h6A;
mem[16'h65AB] = 8'hA5;
mem[16'h65AC] = 8'h6A;
mem[16'h65AD] = 8'h51;
mem[16'h65AE] = 8'h59;
mem[16'h65AF] = 8'h05;
mem[16'h65B0] = 8'h6D;
mem[16'h65B1] = 8'h91;
mem[16'h65B2] = 8'h59;
mem[16'h65B3] = 8'hC8;
mem[16'h65B4] = 8'hA5;
mem[16'h65B5] = 8'h66;
mem[16'h65B6] = 8'h51;
mem[16'h65B7] = 8'h59;
mem[16'h65B8] = 8'h05;
mem[16'h65B9] = 8'h6D;
mem[16'h65BA] = 8'h91;
mem[16'h65BB] = 8'h59;
mem[16'h65BC] = 8'hE6;
mem[16'h65BD] = 8'h56;
mem[16'h65BE] = 8'hE8;
mem[16'h65BF] = 8'hE0;
mem[16'h65C0] = 8'h09;
mem[16'h65C1] = 8'hB0;
mem[16'h65C2] = 8'h03;
mem[16'h65C3] = 8'h4C;
mem[16'h65C4] = 8'h6C;
mem[16'h65C5] = 8'h65;
mem[16'h65C6] = 8'h60;
mem[16'h65C7] = 8'h8D;
mem[16'h65C8] = 8'h88;
mem[16'h65C9] = 8'h65;
mem[16'h65CA] = 8'h8D;
mem[16'h65CB] = 8'h8F;
mem[16'h65CC] = 8'h65;
mem[16'h65CD] = 8'h8C;
mem[16'h65CE] = 8'h89;
mem[16'h65CF] = 8'h65;
mem[16'h65D0] = 8'h8C;
mem[16'h65D1] = 8'h90;
mem[16'h65D2] = 8'h65;
mem[16'h65D3] = 8'h60;
mem[16'h65D4] = 8'h20;
mem[16'h65D5] = 8'h36;
mem[16'h65D6] = 8'h66;
mem[16'h65D7] = 8'hA9;
mem[16'h65D8] = 8'h00;
mem[16'h65D9] = 8'h85;
mem[16'h65DA] = 8'h25;
mem[16'h65DB] = 8'hA9;
mem[16'h65DC] = 8'hF5;
mem[16'h65DD] = 8'h85;
mem[16'h65DE] = 8'h24;
mem[16'h65DF] = 8'hA9;
mem[16'h65E0] = 8'h7D;
mem[16'h65E1] = 8'h85;
mem[16'h65E2] = 8'h59;
mem[16'h65E3] = 8'hA9;
mem[16'h65E4] = 8'h66;
mem[16'h65E5] = 8'h85;
mem[16'h65E6] = 8'h5A;
mem[16'h65E7] = 8'h20;
mem[16'h65E8] = 8'hD5;
mem[16'h65E9] = 8'h67;
mem[16'h65EA] = 8'hA9;
mem[16'h65EB] = 8'h00;
mem[16'h65EC] = 8'h85;
mem[16'h65ED] = 8'h25;
mem[16'h65EE] = 8'hA9;
mem[16'h65EF] = 8'h01;
mem[16'h65F0] = 8'h85;
mem[16'h65F1] = 8'h24;
mem[16'h65F2] = 8'hAD;
mem[16'h65F3] = 8'hD4;
mem[16'h65F4] = 8'h67;
mem[16'h65F5] = 8'hF0;
mem[16'h65F6] = 8'h03;
mem[16'h65F7] = 8'h20;
mem[16'h65F8] = 8'hDA;
mem[16'h65F9] = 8'hFD;
mem[16'h65FA] = 8'hAD;
mem[16'h65FB] = 8'hD3;
mem[16'h65FC] = 8'h67;
mem[16'h65FD] = 8'h20;
mem[16'h65FE] = 8'hDA;
mem[16'h65FF] = 8'hFD;
mem[16'h6600] = 8'hAD;
mem[16'h6601] = 8'hD2;
mem[16'h6602] = 8'h67;
mem[16'h6603] = 8'h20;
mem[16'h6604] = 8'hDA;
mem[16'h6605] = 8'hFD;
mem[16'h6606] = 8'hA9;
mem[16'h6607] = 8'h00;
mem[16'h6608] = 8'h85;
mem[16'h6609] = 8'h25;
mem[16'h660A] = 8'hA9;
mem[16'h660B] = 8'hF7;
mem[16'h660C] = 8'h85;
mem[16'h660D] = 8'h24;
mem[16'h660E] = 8'hA9;
mem[16'h660F] = 8'h73;
mem[16'h6610] = 8'h85;
mem[16'h6611] = 8'h59;
mem[16'h6612] = 8'hA9;
mem[16'h6613] = 8'h66;
mem[16'h6614] = 8'h85;
mem[16'h6615] = 8'h5A;
mem[16'h6616] = 8'h20;
mem[16'h6617] = 8'hD5;
mem[16'h6618] = 8'h67;
mem[16'h6619] = 8'hA9;
mem[16'h661A] = 8'h00;
mem[16'h661B] = 8'h85;
mem[16'h661C] = 8'h25;
mem[16'h661D] = 8'hA9;
mem[16'h661E] = 8'h01;
mem[16'h661F] = 8'h85;
mem[16'h6620] = 8'h24;
mem[16'h6621] = 8'hAD;
mem[16'h6622] = 8'h6F;
mem[16'h6623] = 8'h66;
mem[16'h6624] = 8'hF0;
mem[16'h6625] = 8'h03;
mem[16'h6626] = 8'h20;
mem[16'h6627] = 8'hDA;
mem[16'h6628] = 8'hFD;
mem[16'h6629] = 8'hAD;
mem[16'h662A] = 8'h6E;
mem[16'h662B] = 8'h66;
mem[16'h662C] = 8'h20;
mem[16'h662D] = 8'hDA;
mem[16'h662E] = 8'hFD;
mem[16'h662F] = 8'hAD;
mem[16'h6630] = 8'h6D;
mem[16'h6631] = 8'h66;
mem[16'h6632] = 8'h20;
mem[16'h6633] = 8'hDA;
mem[16'h6634] = 8'hFD;
mem[16'h6635] = 8'h60;
mem[16'h6636] = 8'hAD;
mem[16'h6637] = 8'hD4;
mem[16'h6638] = 8'h67;
mem[16'h6639] = 8'hCD;
mem[16'h663A] = 8'h6F;
mem[16'h663B] = 8'h66;
mem[16'h663C] = 8'h90;
mem[16'h663D] = 8'h2E;
mem[16'h663E] = 8'hF0;
mem[16'h663F] = 8'h03;
mem[16'h6640] = 8'h4C;
mem[16'h6641] = 8'h5A;
mem[16'h6642] = 8'h66;
mem[16'h6643] = 8'hAD;
mem[16'h6644] = 8'hD3;
mem[16'h6645] = 8'h67;
mem[16'h6646] = 8'hCD;
mem[16'h6647] = 8'h6E;
mem[16'h6648] = 8'h66;
mem[16'h6649] = 8'h90;
mem[16'h664A] = 8'h21;
mem[16'h664B] = 8'hF0;
mem[16'h664C] = 8'h03;
mem[16'h664D] = 8'h4C;
mem[16'h664E] = 8'h5A;
mem[16'h664F] = 8'h66;
mem[16'h6650] = 8'hAD;
mem[16'h6651] = 8'hD2;
mem[16'h6652] = 8'h67;
mem[16'h6653] = 8'hCD;
mem[16'h6654] = 8'h6D;
mem[16'h6655] = 8'h66;
mem[16'h6656] = 8'h90;
mem[16'h6657] = 8'h14;
mem[16'h6658] = 8'hF0;
mem[16'h6659] = 8'h12;
mem[16'h665A] = 8'hAD;
mem[16'h665B] = 8'hD2;
mem[16'h665C] = 8'h67;
mem[16'h665D] = 8'h8D;
mem[16'h665E] = 8'h6D;
mem[16'h665F] = 8'h66;
mem[16'h6660] = 8'hAD;
mem[16'h6661] = 8'hD3;
mem[16'h6662] = 8'h67;
mem[16'h6663] = 8'h8D;
mem[16'h6664] = 8'h6E;
mem[16'h6665] = 8'h66;
mem[16'h6666] = 8'hAD;
mem[16'h6667] = 8'hD4;
mem[16'h6668] = 8'h67;
mem[16'h6669] = 8'h8D;
mem[16'h666A] = 8'h6F;
mem[16'h666B] = 8'h66;
mem[16'h666C] = 8'h60;
mem[16'h666D] = 8'h00;
mem[16'h666E] = 8'h00;
mem[16'h666F] = 8'h00;
mem[16'h6670] = 8'h00;
mem[16'h6671] = 8'h00;
mem[16'h6672] = 8'h00;
mem[16'h6673] = 8'hA0;
mem[16'h6674] = 8'hC8;
mem[16'h6675] = 8'hE9;
mem[16'h6676] = 8'hA0;
mem[16'h6677] = 8'hD3;
mem[16'h6678] = 8'hE3;
mem[16'h6679] = 8'hEF;
mem[16'h667A] = 8'hF2;
mem[16'h667B] = 8'hE5;
mem[16'h667C] = 8'h00;
mem[16'h667D] = 8'hA0;
mem[16'h667E] = 8'hD9;
mem[16'h667F] = 8'hEF;
mem[16'h6680] = 8'hF5;
mem[16'h6681] = 8'hF2;
mem[16'h6682] = 8'hA0;
mem[16'h6683] = 8'hD3;
mem[16'h6684] = 8'hE3;
mem[16'h6685] = 8'hEF;
mem[16'h6686] = 8'hF2;
mem[16'h6687] = 8'hE5;
mem[16'h6688] = 8'h00;
mem[16'h6689] = 8'hF8;
mem[16'h668A] = 8'h18;
mem[16'h668B] = 8'h6D;
mem[16'h668C] = 8'hD2;
mem[16'h668D] = 8'h67;
mem[16'h668E] = 8'h8D;
mem[16'h668F] = 8'hD2;
mem[16'h6690] = 8'h67;
mem[16'h6691] = 8'h90;
mem[16'h6692] = 8'h12;
mem[16'h6693] = 8'hAD;
mem[16'h6694] = 8'hD3;
mem[16'h6695] = 8'h67;
mem[16'h6696] = 8'h69;
mem[16'h6697] = 8'h00;
mem[16'h6698] = 8'h8D;
mem[16'h6699] = 8'hD3;
mem[16'h669A] = 8'h67;
mem[16'h669B] = 8'h90;
mem[16'h669C] = 8'h08;
mem[16'h669D] = 8'hAD;
mem[16'h669E] = 8'hD4;
mem[16'h669F] = 8'h67;
mem[16'h66A0] = 8'h69;
mem[16'h66A1] = 8'h00;
mem[16'h66A2] = 8'h8D;
mem[16'h66A3] = 8'hD4;
mem[16'h66A4] = 8'h67;
mem[16'h66A5] = 8'hD8;
mem[16'h66A6] = 8'h20;
mem[16'h66A7] = 8'h36;
mem[16'h66A8] = 8'h66;
mem[16'h66A9] = 8'h20;
mem[16'h66AA] = 8'hB5;
mem[16'h66AB] = 8'h66;
mem[16'h66AC] = 8'h60;
mem[16'h66AD] = 8'hF8;
mem[16'h66AE] = 8'h18;
mem[16'h66AF] = 8'h6D;
mem[16'h66B0] = 8'hD3;
mem[16'h66B1] = 8'h67;
mem[16'h66B2] = 8'h4C;
mem[16'h66B3] = 8'h98;
mem[16'h66B4] = 8'h66;
mem[16'h66B5] = 8'hA9;
mem[16'h66B6] = 8'h00;
mem[16'h66B7] = 8'h85;
mem[16'h66B8] = 8'h25;
mem[16'h66B9] = 8'hA9;
mem[16'h66BA] = 8'h1F;
mem[16'h66BB] = 8'h85;
mem[16'h66BC] = 8'h24;
mem[16'h66BD] = 8'hAD;
mem[16'h66BE] = 8'hD1;
mem[16'h66BF] = 8'h67;
mem[16'h66C0] = 8'hCD;
mem[16'h66C1] = 8'hD4;
mem[16'h66C2] = 8'h67;
mem[16'h66C3] = 8'hF0;
mem[16'h66C4] = 8'h10;
mem[16'h66C5] = 8'h20;
mem[16'h66C6] = 8'hDA;
mem[16'h66C7] = 8'hFD;
mem[16'h66C8] = 8'hA2;
mem[16'h66C9] = 8'h1F;
mem[16'h66CA] = 8'h86;
mem[16'h66CB] = 8'h24;
mem[16'h66CC] = 8'hAD;
mem[16'h66CD] = 8'hD4;
mem[16'h66CE] = 8'h67;
mem[16'h66CF] = 8'h8D;
mem[16'h66D0] = 8'hD1;
mem[16'h66D1] = 8'h67;
mem[16'h66D2] = 8'h20;
mem[16'h66D3] = 8'hDA;
mem[16'h66D4] = 8'hFD;
mem[16'h66D5] = 8'hAD;
mem[16'h66D6] = 8'hD0;
mem[16'h66D7] = 8'h67;
mem[16'h66D8] = 8'hCD;
mem[16'h66D9] = 8'hD3;
mem[16'h66DA] = 8'h67;
mem[16'h66DB] = 8'hF0;
mem[16'h66DC] = 8'h14;
mem[16'h66DD] = 8'hA2;
mem[16'h66DE] = 8'h21;
mem[16'h66DF] = 8'h86;
mem[16'h66E0] = 8'h24;
mem[16'h66E1] = 8'h20;
mem[16'h66E2] = 8'hDA;
mem[16'h66E3] = 8'hFD;
mem[16'h66E4] = 8'hA2;
mem[16'h66E5] = 8'h21;
mem[16'h66E6] = 8'h86;
mem[16'h66E7] = 8'h24;
mem[16'h66E8] = 8'hAD;
mem[16'h66E9] = 8'hD3;
mem[16'h66EA] = 8'h67;
mem[16'h66EB] = 8'h8D;
mem[16'h66EC] = 8'hD0;
mem[16'h66ED] = 8'h67;
mem[16'h66EE] = 8'h20;
mem[16'h66EF] = 8'hDA;
mem[16'h66F0] = 8'hFD;
mem[16'h66F1] = 8'hAD;
mem[16'h66F2] = 8'hCF;
mem[16'h66F3] = 8'h67;
mem[16'h66F4] = 8'hCD;
mem[16'h66F5] = 8'hD2;
mem[16'h66F6] = 8'h67;
mem[16'h66F7] = 8'hF0;
mem[16'h66F8] = 8'h14;
mem[16'h66F9] = 8'hA2;
mem[16'h66FA] = 8'h23;
mem[16'h66FB] = 8'h86;
mem[16'h66FC] = 8'h24;
mem[16'h66FD] = 8'h20;
mem[16'h66FE] = 8'hDA;
mem[16'h66FF] = 8'hFD;
mem[16'h6700] = 8'hA2;
mem[16'h6701] = 8'h23;
mem[16'h6702] = 8'h86;
mem[16'h6703] = 8'h24;
mem[16'h6704] = 8'hAD;
mem[16'h6705] = 8'hD2;
mem[16'h6706] = 8'h67;
mem[16'h6707] = 8'h8D;
mem[16'h6708] = 8'hCF;
mem[16'h6709] = 8'h67;
mem[16'h670A] = 8'h20;
mem[16'h670B] = 8'hDA;
mem[16'h670C] = 8'hFD;
mem[16'h670D] = 8'hA9;
mem[16'h670E] = 8'h0A;
mem[16'h670F] = 8'h85;
mem[16'h6710] = 8'h24;
mem[16'h6711] = 8'hAD;
mem[16'h6712] = 8'h72;
mem[16'h6713] = 8'h66;
mem[16'h6714] = 8'hCD;
mem[16'h6715] = 8'h6F;
mem[16'h6716] = 8'h66;
mem[16'h6717] = 8'hF0;
mem[16'h6718] = 8'h10;
mem[16'h6719] = 8'h20;
mem[16'h671A] = 8'hDA;
mem[16'h671B] = 8'hFD;
mem[16'h671C] = 8'hA2;
mem[16'h671D] = 8'h0A;
mem[16'h671E] = 8'h86;
mem[16'h671F] = 8'h24;
mem[16'h6720] = 8'hAD;
mem[16'h6721] = 8'h6F;
mem[16'h6722] = 8'h66;
mem[16'h6723] = 8'h8D;
mem[16'h6724] = 8'h72;
mem[16'h6725] = 8'h66;
mem[16'h6726] = 8'h20;
mem[16'h6727] = 8'hDA;
mem[16'h6728] = 8'hFD;
mem[16'h6729] = 8'hAD;
mem[16'h672A] = 8'h71;
mem[16'h672B] = 8'h66;
mem[16'h672C] = 8'hCD;
mem[16'h672D] = 8'h6E;
mem[16'h672E] = 8'h66;
mem[16'h672F] = 8'hF0;
mem[16'h6730] = 8'h14;
mem[16'h6731] = 8'hA2;
mem[16'h6732] = 8'h0C;
mem[16'h6733] = 8'h86;
mem[16'h6734] = 8'h24;
mem[16'h6735] = 8'h20;
mem[16'h6736] = 8'hDA;
mem[16'h6737] = 8'hFD;
mem[16'h6738] = 8'hA2;
mem[16'h6739] = 8'h0C;
mem[16'h673A] = 8'h86;
mem[16'h673B] = 8'h24;
mem[16'h673C] = 8'hAD;
mem[16'h673D] = 8'h6E;
mem[16'h673E] = 8'h66;
mem[16'h673F] = 8'h8D;
mem[16'h6740] = 8'h71;
mem[16'h6741] = 8'h66;
mem[16'h6742] = 8'h20;
mem[16'h6743] = 8'hDA;
mem[16'h6744] = 8'hFD;
mem[16'h6745] = 8'hAD;
mem[16'h6746] = 8'h70;
mem[16'h6747] = 8'h66;
mem[16'h6748] = 8'hCD;
mem[16'h6749] = 8'h6D;
mem[16'h674A] = 8'h66;
mem[16'h674B] = 8'hF0;
mem[16'h674C] = 8'h14;
mem[16'h674D] = 8'hA2;
mem[16'h674E] = 8'h0E;
mem[16'h674F] = 8'h86;
mem[16'h6750] = 8'h24;
mem[16'h6751] = 8'h20;
mem[16'h6752] = 8'hDA;
mem[16'h6753] = 8'hFD;
mem[16'h6754] = 8'hA2;
mem[16'h6755] = 8'h0E;
mem[16'h6756] = 8'h86;
mem[16'h6757] = 8'h24;
mem[16'h6758] = 8'hAD;
mem[16'h6759] = 8'h6D;
mem[16'h675A] = 8'h66;
mem[16'h675B] = 8'h8D;
mem[16'h675C] = 8'h70;
mem[16'h675D] = 8'h66;
mem[16'h675E] = 8'h20;
mem[16'h675F] = 8'hDA;
mem[16'h6760] = 8'hFD;
mem[16'h6761] = 8'h60;
mem[16'h6762] = 8'hA9;
mem[16'h6763] = 8'h00;
mem[16'h6764] = 8'h85;
mem[16'h6765] = 8'h25;
mem[16'h6766] = 8'hA9;
mem[16'h6767] = 8'h00;
mem[16'h6768] = 8'h85;
mem[16'h6769] = 8'h24;
mem[16'h676A] = 8'hA9;
mem[16'h676B] = 8'h73;
mem[16'h676C] = 8'h85;
mem[16'h676D] = 8'h59;
mem[16'h676E] = 8'hA9;
mem[16'h676F] = 8'h66;
mem[16'h6770] = 8'h85;
mem[16'h6771] = 8'h5A;
mem[16'h6772] = 8'h20;
mem[16'h6773] = 8'hD5;
mem[16'h6774] = 8'h67;
mem[16'h6775] = 8'hA9;
mem[16'h6776] = 8'h00;
mem[16'h6777] = 8'h85;
mem[16'h6778] = 8'h25;
mem[16'h6779] = 8'hA9;
mem[16'h677A] = 8'h13;
mem[16'h677B] = 8'h85;
mem[16'h677C] = 8'h24;
mem[16'h677D] = 8'hA9;
mem[16'h677E] = 8'h7D;
mem[16'h677F] = 8'h85;
mem[16'h6780] = 8'h59;
mem[16'h6781] = 8'hA9;
mem[16'h6782] = 8'h66;
mem[16'h6783] = 8'h85;
mem[16'h6784] = 8'h5A;
mem[16'h6785] = 8'h20;
mem[16'h6786] = 8'hD5;
mem[16'h6787] = 8'h67;
mem[16'h6788] = 8'hA9;
mem[16'h6789] = 8'h00;
mem[16'h678A] = 8'h85;
mem[16'h678B] = 8'h25;
mem[16'h678C] = 8'hA9;
mem[16'h678D] = 8'h1F;
mem[16'h678E] = 8'h85;
mem[16'h678F] = 8'h24;
mem[16'h6790] = 8'hAD;
mem[16'h6791] = 8'hD4;
mem[16'h6792] = 8'h67;
mem[16'h6793] = 8'h8D;
mem[16'h6794] = 8'hD1;
mem[16'h6795] = 8'h67;
mem[16'h6796] = 8'h20;
mem[16'h6797] = 8'hDA;
mem[16'h6798] = 8'hFD;
mem[16'h6799] = 8'hAD;
mem[16'h679A] = 8'hD3;
mem[16'h679B] = 8'h67;
mem[16'h679C] = 8'h8D;
mem[16'h679D] = 8'hD0;
mem[16'h679E] = 8'h67;
mem[16'h679F] = 8'h20;
mem[16'h67A0] = 8'hDA;
mem[16'h67A1] = 8'hFD;
mem[16'h67A2] = 8'hAD;
mem[16'h67A3] = 8'hD2;
mem[16'h67A4] = 8'h67;
mem[16'h67A5] = 8'h8D;
mem[16'h67A6] = 8'hCF;
mem[16'h67A7] = 8'h67;
mem[16'h67A8] = 8'h20;
mem[16'h67A9] = 8'hDA;
mem[16'h67AA] = 8'hFD;
mem[16'h67AB] = 8'hA9;
mem[16'h67AC] = 8'h00;
mem[16'h67AD] = 8'h85;
mem[16'h67AE] = 8'h25;
mem[16'h67AF] = 8'hA9;
mem[16'h67B0] = 8'h0A;
mem[16'h67B1] = 8'h85;
mem[16'h67B2] = 8'h24;
mem[16'h67B3] = 8'hAD;
mem[16'h67B4] = 8'h6F;
mem[16'h67B5] = 8'h66;
mem[16'h67B6] = 8'h8D;
mem[16'h67B7] = 8'h72;
mem[16'h67B8] = 8'h66;
mem[16'h67B9] = 8'h20;
mem[16'h67BA] = 8'hDA;
mem[16'h67BB] = 8'hFD;
mem[16'h67BC] = 8'hAD;
mem[16'h67BD] = 8'h6E;
mem[16'h67BE] = 8'h66;
mem[16'h67BF] = 8'h8D;
mem[16'h67C0] = 8'h71;
mem[16'h67C1] = 8'h66;
mem[16'h67C2] = 8'h20;
mem[16'h67C3] = 8'hDA;
mem[16'h67C4] = 8'hFD;
mem[16'h67C5] = 8'hAD;
mem[16'h67C6] = 8'h6D;
mem[16'h67C7] = 8'h66;
mem[16'h67C8] = 8'h8D;
mem[16'h67C9] = 8'h70;
mem[16'h67CA] = 8'h66;
mem[16'h67CB] = 8'h20;
mem[16'h67CC] = 8'hDA;
mem[16'h67CD] = 8'hFD;
mem[16'h67CE] = 8'h60;
mem[16'h67CF] = 8'h00;
mem[16'h67D0] = 8'h00;
mem[16'h67D1] = 8'h00;
mem[16'h67D2] = 8'h00;
mem[16'h67D3] = 8'h00;
mem[16'h67D4] = 8'h00;
mem[16'h67D5] = 8'hA0;
mem[16'h67D6] = 8'h00;
mem[16'h67D7] = 8'hB1;
mem[16'h67D8] = 8'h59;
mem[16'h67D9] = 8'hF0;
mem[16'h67DA] = 8'h07;
mem[16'h67DB] = 8'h20;
mem[16'h67DC] = 8'hED;
mem[16'h67DD] = 8'hFD;
mem[16'h67DE] = 8'hC8;
mem[16'h67DF] = 8'h4C;
mem[16'h67E0] = 8'hD7;
mem[16'h67E1] = 8'h67;
mem[16'h67E2] = 8'h20;
mem[16'h67E3] = 8'h8E;
mem[16'h67E4] = 8'hFD;
mem[16'h67E5] = 8'h60;
mem[16'h67E6] = 8'hA2;
mem[16'h67E7] = 8'h00;
mem[16'h67E8] = 8'hA4;
mem[16'h67E9] = 8'h56;
mem[16'h67EA] = 8'hB9;
mem[16'h67EB] = 8'hD5;
mem[16'h67EC] = 8'h8E;
mem[16'h67ED] = 8'h85;
mem[16'h67EE] = 8'h59;
mem[16'h67EF] = 8'hB9;
mem[16'h67F0] = 8'h95;
mem[16'h67F1] = 8'h8F;
mem[16'h67F2] = 8'h45;
mem[16'h67F3] = 8'h64;
mem[16'h67F4] = 8'h85;
mem[16'h67F5] = 8'h5A;
mem[16'h67F6] = 8'hA4;
mem[16'h67F7] = 8'h57;
mem[16'h67F8] = 8'hB9;
mem[16'h67F9] = 8'h3E;
mem[16'h67FA] = 8'h8C;
mem[16'h67FB] = 8'h85;
mem[16'h67FC] = 8'h5C;
mem[16'h67FD] = 8'hB9;
mem[16'h67FE] = 8'h56;
mem[16'h67FF] = 8'h8D;
mem[16'h6800] = 8'hA8;
mem[16'h6801] = 8'hBD;
mem[16'h6802] = 8'h2F;
mem[16'h6803] = 8'h60;
mem[16'h6804] = 8'h29;
mem[16'h6805] = 8'h80;
mem[16'h6806] = 8'h85;
mem[16'h6807] = 8'h6D;
mem[16'h6808] = 8'hBD;
mem[16'h6809] = 8'h2F;
mem[16'h680A] = 8'h60;
mem[16'h680B] = 8'h29;
mem[16'h680C] = 8'h7F;
mem[16'h680D] = 8'h85;
mem[16'h680E] = 8'h66;
mem[16'h680F] = 8'hE8;
mem[16'h6810] = 8'hBD;
mem[16'h6811] = 8'h2F;
mem[16'h6812] = 8'h60;
mem[16'h6813] = 8'h29;
mem[16'h6814] = 8'h7F;
mem[16'h6815] = 8'h85;
mem[16'h6816] = 8'h67;
mem[16'h6817] = 8'hE8;
mem[16'h6818] = 8'hBD;
mem[16'h6819] = 8'h2F;
mem[16'h681A] = 8'h60;
mem[16'h681B] = 8'h29;
mem[16'h681C] = 8'h7F;
mem[16'h681D] = 8'h85;
mem[16'h681E] = 8'h68;
mem[16'h681F] = 8'hA9;
mem[16'h6820] = 8'h00;
mem[16'h6821] = 8'h85;
mem[16'h6822] = 8'h6B;
mem[16'h6823] = 8'h85;
mem[16'h6824] = 8'h6C;
mem[16'h6825] = 8'h85;
mem[16'h6826] = 8'h6A;
mem[16'h6827] = 8'h85;
mem[16'h6828] = 8'h69;
mem[16'h6829] = 8'hA5;
mem[16'h682A] = 8'h5C;
mem[16'h682B] = 8'hC9;
mem[16'h682C] = 8'h01;
mem[16'h682D] = 8'hF0;
mem[16'h682E] = 8'h29;
mem[16'h682F] = 8'h46;
mem[16'h6830] = 8'h67;
mem[16'h6831] = 8'h66;
mem[16'h6832] = 8'h6B;
mem[16'h6833] = 8'h46;
mem[16'h6834] = 8'h66;
mem[16'h6835] = 8'h66;
mem[16'h6836] = 8'h6A;
mem[16'h6837] = 8'h46;
mem[16'h6838] = 8'h68;
mem[16'h6839] = 8'h66;
mem[16'h683A] = 8'h6C;
mem[16'h683B] = 8'h06;
mem[16'h683C] = 8'h5C;
mem[16'h683D] = 8'h24;
mem[16'h683E] = 8'h5C;
mem[16'h683F] = 8'h10;
mem[16'h6840] = 8'hEE;
mem[16'h6841] = 8'hA5;
mem[16'h6842] = 8'h68;
mem[16'h6843] = 8'h85;
mem[16'h6844] = 8'h69;
mem[16'h6845] = 8'hA5;
mem[16'h6846] = 8'h6C;
mem[16'h6847] = 8'h4A;
mem[16'h6848] = 8'h05;
mem[16'h6849] = 8'h67;
mem[16'h684A] = 8'h85;
mem[16'h684B] = 8'h68;
mem[16'h684C] = 8'hA5;
mem[16'h684D] = 8'h6B;
mem[16'h684E] = 8'h4A;
mem[16'h684F] = 8'h05;
mem[16'h6850] = 8'h66;
mem[16'h6851] = 8'h85;
mem[16'h6852] = 8'h67;
mem[16'h6853] = 8'hA5;
mem[16'h6854] = 8'h6A;
mem[16'h6855] = 8'h4A;
mem[16'h6856] = 8'h85;
mem[16'h6857] = 8'h66;
mem[16'h6858] = 8'hA5;
mem[16'h6859] = 8'h66;
mem[16'h685A] = 8'h05;
mem[16'h685B] = 8'h6D;
mem[16'h685C] = 8'h51;
mem[16'h685D] = 8'h59;
mem[16'h685E] = 8'h91;
mem[16'h685F] = 8'h59;
mem[16'h6860] = 8'hC8;
mem[16'h6861] = 8'hA5;
mem[16'h6862] = 8'h67;
mem[16'h6863] = 8'h05;
mem[16'h6864] = 8'h6D;
mem[16'h6865] = 8'h51;
mem[16'h6866] = 8'h59;
mem[16'h6867] = 8'h91;
mem[16'h6868] = 8'h59;
mem[16'h6869] = 8'hC8;
mem[16'h686A] = 8'hA5;
mem[16'h686B] = 8'h68;
mem[16'h686C] = 8'h05;
mem[16'h686D] = 8'h6D;
mem[16'h686E] = 8'h51;
mem[16'h686F] = 8'h59;
mem[16'h6870] = 8'h91;
mem[16'h6871] = 8'h59;
mem[16'h6872] = 8'hC8;
mem[16'h6873] = 8'hA5;
mem[16'h6874] = 8'h69;
mem[16'h6875] = 8'h05;
mem[16'h6876] = 8'h6D;
mem[16'h6877] = 8'h51;
mem[16'h6878] = 8'h59;
mem[16'h6879] = 8'h91;
mem[16'h687A] = 8'h59;
mem[16'h687B] = 8'hE6;
mem[16'h687C] = 8'h56;
mem[16'h687D] = 8'hE8;
mem[16'h687E] = 8'hE0;
mem[16'h687F] = 8'h18;
mem[16'h6880] = 8'hF0;
mem[16'h6881] = 8'h03;
mem[16'h6882] = 8'h4C;
mem[16'h6883] = 8'hE8;
mem[16'h6884] = 8'h67;
mem[16'h6885] = 8'h60;
mem[16'h6886] = 8'h8D;
mem[16'h6887] = 8'h02;
mem[16'h6888] = 8'h68;
mem[16'h6889] = 8'h8D;
mem[16'h688A] = 8'h09;
mem[16'h688B] = 8'h68;
mem[16'h688C] = 8'h8D;
mem[16'h688D] = 8'h11;
mem[16'h688E] = 8'h68;
mem[16'h688F] = 8'h8D;
mem[16'h6890] = 8'h19;
mem[16'h6891] = 8'h68;
mem[16'h6892] = 8'h8C;
mem[16'h6893] = 8'h03;
mem[16'h6894] = 8'h68;
mem[16'h6895] = 8'h8C;
mem[16'h6896] = 8'h0A;
mem[16'h6897] = 8'h68;
mem[16'h6898] = 8'h8C;
mem[16'h6899] = 8'h12;
mem[16'h689A] = 8'h68;
mem[16'h689B] = 8'h8C;
mem[16'h689C] = 8'h1A;
mem[16'h689D] = 8'h68;
mem[16'h689E] = 8'h60;
mem[16'h689F] = 8'hA2;
mem[16'h68A0] = 8'h00;
mem[16'h68A1] = 8'hA4;
mem[16'h68A2] = 8'h56;
mem[16'h68A3] = 8'hC0;
mem[16'h68A4] = 8'hC0;
mem[16'h68A5] = 8'h90;
mem[16'h68A6] = 8'h06;
mem[16'h68A7] = 8'h20;
mem[16'h68A8] = 8'hDD;
mem[16'h68A9] = 8'hFB;
mem[16'h68AA] = 8'h4C;
mem[16'h68AB] = 8'h0D;
mem[16'h68AC] = 8'h69;
mem[16'h68AD] = 8'hB9;
mem[16'h68AE] = 8'hD5;
mem[16'h68AF] = 8'h8E;
mem[16'h68B0] = 8'h85;
mem[16'h68B1] = 8'h59;
mem[16'h68B2] = 8'hB9;
mem[16'h68B3] = 8'h95;
mem[16'h68B4] = 8'h8F;
mem[16'h68B5] = 8'h85;
mem[16'h68B6] = 8'h5A;
mem[16'h68B7] = 8'hA4;
mem[16'h68B8] = 8'h57;
mem[16'h68B9] = 8'hB9;
mem[16'h68BA] = 8'h56;
mem[16'h68BB] = 8'h8D;
mem[16'h68BC] = 8'hA8;
mem[16'h68BD] = 8'hBD;
mem[16'h68BE] = 8'h00;
mem[16'h68BF] = 8'h00;
mem[16'h68C0] = 8'h29;
mem[16'h68C1] = 8'h80;
mem[16'h68C2] = 8'h85;
mem[16'h68C3] = 8'h6D;
mem[16'h68C4] = 8'hBD;
mem[16'h68C5] = 8'h00;
mem[16'h68C6] = 8'h00;
mem[16'h68C7] = 8'h29;
mem[16'h68C8] = 8'h7F;
mem[16'h68C9] = 8'h51;
mem[16'h68CA] = 8'h59;
mem[16'h68CB] = 8'h05;
mem[16'h68CC] = 8'h6D;
mem[16'h68CD] = 8'h91;
mem[16'h68CE] = 8'h59;
mem[16'h68CF] = 8'hE8;
mem[16'h68D0] = 8'hC8;
mem[16'h68D1] = 8'hBD;
mem[16'h68D2] = 8'h00;
mem[16'h68D3] = 8'h00;
mem[16'h68D4] = 8'h29;
mem[16'h68D5] = 8'h7F;
mem[16'h68D6] = 8'h51;
mem[16'h68D7] = 8'h59;
mem[16'h68D8] = 8'h05;
mem[16'h68D9] = 8'h6D;
mem[16'h68DA] = 8'h91;
mem[16'h68DB] = 8'h59;
mem[16'h68DC] = 8'hC8;
mem[16'h68DD] = 8'hE8;
mem[16'h68DE] = 8'hBD;
mem[16'h68DF] = 8'h00;
mem[16'h68E0] = 8'h00;
mem[16'h68E1] = 8'h29;
mem[16'h68E2] = 8'h7F;
mem[16'h68E3] = 8'h51;
mem[16'h68E4] = 8'h59;
mem[16'h68E5] = 8'h05;
mem[16'h68E6] = 8'h6D;
mem[16'h68E7] = 8'h91;
mem[16'h68E8] = 8'h59;
mem[16'h68E9] = 8'hC8;
mem[16'h68EA] = 8'hE8;
mem[16'h68EB] = 8'hBD;
mem[16'h68EC] = 8'h00;
mem[16'h68ED] = 8'h00;
mem[16'h68EE] = 8'h29;
mem[16'h68EF] = 8'h7F;
mem[16'h68F0] = 8'h51;
mem[16'h68F1] = 8'h59;
mem[16'h68F2] = 8'h05;
mem[16'h68F3] = 8'h6D;
mem[16'h68F4] = 8'h91;
mem[16'h68F5] = 8'h59;
mem[16'h68F6] = 8'hC8;
mem[16'h68F7] = 8'hE8;
mem[16'h68F8] = 8'hBD;
mem[16'h68F9] = 8'h00;
mem[16'h68FA] = 8'h00;
mem[16'h68FB] = 8'h29;
mem[16'h68FC] = 8'h7F;
mem[16'h68FD] = 8'h51;
mem[16'h68FE] = 8'h59;
mem[16'h68FF] = 8'h05;
mem[16'h6900] = 8'h6D;
mem[16'h6901] = 8'h91;
mem[16'h6902] = 8'h59;
mem[16'h6903] = 8'hE6;
mem[16'h6904] = 8'h56;
mem[16'h6905] = 8'hE8;
mem[16'h6906] = 8'hE0;
mem[16'h6907] = 8'h1E;
mem[16'h6908] = 8'hB0;
mem[16'h6909] = 8'h03;
mem[16'h690A] = 8'h4C;
mem[16'h690B] = 8'hA1;
mem[16'h690C] = 8'h68;
mem[16'h690D] = 8'h60;
mem[16'h690E] = 8'h8D;
mem[16'h690F] = 8'hBE;
mem[16'h6910] = 8'h68;
mem[16'h6911] = 8'h8D;
mem[16'h6912] = 8'hC5;
mem[16'h6913] = 8'h68;
mem[16'h6914] = 8'h8D;
mem[16'h6915] = 8'hD2;
mem[16'h6916] = 8'h68;
mem[16'h6917] = 8'h8D;
mem[16'h6918] = 8'hDF;
mem[16'h6919] = 8'h68;
mem[16'h691A] = 8'h8D;
mem[16'h691B] = 8'hEC;
mem[16'h691C] = 8'h68;
mem[16'h691D] = 8'h8D;
mem[16'h691E] = 8'hF9;
mem[16'h691F] = 8'h68;
mem[16'h6920] = 8'h8C;
mem[16'h6921] = 8'hBF;
mem[16'h6922] = 8'h68;
mem[16'h6923] = 8'h8C;
mem[16'h6924] = 8'hC6;
mem[16'h6925] = 8'h68;
mem[16'h6926] = 8'h8C;
mem[16'h6927] = 8'hD3;
mem[16'h6928] = 8'h68;
mem[16'h6929] = 8'h8C;
mem[16'h692A] = 8'hE0;
mem[16'h692B] = 8'h68;
mem[16'h692C] = 8'h8C;
mem[16'h692D] = 8'hED;
mem[16'h692E] = 8'h68;
mem[16'h692F] = 8'h8C;
mem[16'h6930] = 8'hFA;
mem[16'h6931] = 8'h68;
mem[16'h6932] = 8'h60;
mem[16'h6933] = 8'hA2;
mem[16'h6934] = 8'h00;
mem[16'h6935] = 8'h86;
mem[16'h6936] = 8'h76;
mem[16'h6937] = 8'hA4;
mem[16'h6938] = 8'h56;
mem[16'h6939] = 8'hC0;
mem[16'h693A] = 8'hC0;
mem[16'h693B] = 8'h90;
mem[16'h693C] = 8'h06;
mem[16'h693D] = 8'h20;
mem[16'h693E] = 8'hDD;
mem[16'h693F] = 8'hFB;
mem[16'h6940] = 8'h4C;
mem[16'h6941] = 8'hFF;
mem[16'h6942] = 8'h69;
mem[16'h6943] = 8'hB9;
mem[16'h6944] = 8'hD5;
mem[16'h6945] = 8'h8E;
mem[16'h6946] = 8'h85;
mem[16'h6947] = 8'h59;
mem[16'h6948] = 8'hB9;
mem[16'h6949] = 8'h95;
mem[16'h694A] = 8'h8F;
mem[16'h694B] = 8'h85;
mem[16'h694C] = 8'h5A;
mem[16'h694D] = 8'hA4;
mem[16'h694E] = 8'h57;
mem[16'h694F] = 8'hB9;
mem[16'h6950] = 8'h3E;
mem[16'h6951] = 8'h8C;
mem[16'h6952] = 8'h85;
mem[16'h6953] = 8'h5C;
mem[16'h6954] = 8'hB9;
mem[16'h6955] = 8'h56;
mem[16'h6956] = 8'h8D;
mem[16'h6957] = 8'hA8;
mem[16'h6958] = 8'hBD;
mem[16'h6959] = 8'hF3;
mem[16'h695A] = 8'h4C;
mem[16'h695B] = 8'h29;
mem[16'h695C] = 8'h80;
mem[16'h695D] = 8'h85;
mem[16'h695E] = 8'h6D;
mem[16'h695F] = 8'hBD;
mem[16'h6960] = 8'hF3;
mem[16'h6961] = 8'h4C;
mem[16'h6962] = 8'h29;
mem[16'h6963] = 8'h7F;
mem[16'h6964] = 8'h85;
mem[16'h6965] = 8'h66;
mem[16'h6966] = 8'hE8;
mem[16'h6967] = 8'hBD;
mem[16'h6968] = 8'hF3;
mem[16'h6969] = 8'h4C;
mem[16'h696A] = 8'h29;
mem[16'h696B] = 8'h7F;
mem[16'h696C] = 8'h85;
mem[16'h696D] = 8'h67;
mem[16'h696E] = 8'hA9;
mem[16'h696F] = 8'h7F;
mem[16'h6970] = 8'h85;
mem[16'h6971] = 8'h78;
mem[16'h6972] = 8'h85;
mem[16'h6973] = 8'h79;
mem[16'h6974] = 8'hA9;
mem[16'h6975] = 8'h00;
mem[16'h6976] = 8'h85;
mem[16'h6977] = 8'h7A;
mem[16'h6978] = 8'h85;
mem[16'h6979] = 8'h68;
mem[16'h697A] = 8'h46;
mem[16'h697B] = 8'h5C;
mem[16'h697C] = 8'hB0;
mem[16'h697D] = 8'h2A;
mem[16'h697E] = 8'h06;
mem[16'h697F] = 8'h66;
mem[16'h6980] = 8'h06;
mem[16'h6981] = 8'h78;
mem[16'h6982] = 8'h06;
mem[16'h6983] = 8'h66;
mem[16'h6984] = 8'h26;
mem[16'h6985] = 8'h67;
mem[16'h6986] = 8'hA5;
mem[16'h6987] = 8'h67;
mem[16'h6988] = 8'h2A;
mem[16'h6989] = 8'h26;
mem[16'h698A] = 8'h68;
mem[16'h698B] = 8'h06;
mem[16'h698C] = 8'h78;
mem[16'h698D] = 8'h26;
mem[16'h698E] = 8'h79;
mem[16'h698F] = 8'hA5;
mem[16'h6990] = 8'h79;
mem[16'h6991] = 8'h2A;
mem[16'h6992] = 8'h26;
mem[16'h6993] = 8'h7A;
mem[16'h6994] = 8'h46;
mem[16'h6995] = 8'h5C;
mem[16'h6996] = 8'h90;
mem[16'h6997] = 8'hEA;
mem[16'h6998] = 8'h46;
mem[16'h6999] = 8'h66;
mem[16'h699A] = 8'hA5;
mem[16'h699B] = 8'h67;
mem[16'h699C] = 8'h29;
mem[16'h699D] = 8'h7F;
mem[16'h699E] = 8'h85;
mem[16'h699F] = 8'h67;
mem[16'h69A0] = 8'h46;
mem[16'h69A1] = 8'h78;
mem[16'h69A2] = 8'hA5;
mem[16'h69A3] = 8'h79;
mem[16'h69A4] = 8'h29;
mem[16'h69A5] = 8'h7F;
mem[16'h69A6] = 8'h85;
mem[16'h69A7] = 8'h79;
mem[16'h69A8] = 8'h86;
mem[16'h69A9] = 8'h62;
mem[16'h69AA] = 8'hA6;
mem[16'h69AB] = 8'h76;
mem[16'h69AC] = 8'hA5;
mem[16'h69AD] = 8'h77;
mem[16'h69AE] = 8'hD0;
mem[16'h69AF] = 8'h19;
mem[16'h69B0] = 8'hB1;
mem[16'h69B1] = 8'h59;
mem[16'h69B2] = 8'h25;
mem[16'h69B3] = 8'h78;
mem[16'h69B4] = 8'h9D;
mem[16'h69B5] = 8'h06;
mem[16'h69B6] = 8'h6A;
mem[16'h69B7] = 8'hC8;
mem[16'h69B8] = 8'hB1;
mem[16'h69B9] = 8'h59;
mem[16'h69BA] = 8'h25;
mem[16'h69BB] = 8'h79;
mem[16'h69BC] = 8'h9D;
mem[16'h69BD] = 8'h07;
mem[16'h69BE] = 8'h6A;
mem[16'h69BF] = 8'hC8;
mem[16'h69C0] = 8'hB1;
mem[16'h69C1] = 8'h59;
mem[16'h69C2] = 8'h25;
mem[16'h69C3] = 8'h7A;
mem[16'h69C4] = 8'h9D;
mem[16'h69C5] = 8'h08;
mem[16'h69C6] = 8'h6A;
mem[16'h69C7] = 8'h88;
mem[16'h69C8] = 8'h88;
mem[16'h69C9] = 8'hA5;
mem[16'h69CA] = 8'h66;
mem[16'h69CB] = 8'h05;
mem[16'h69CC] = 8'h6D;
mem[16'h69CD] = 8'h51;
mem[16'h69CE] = 8'h59;
mem[16'h69CF] = 8'h5D;
mem[16'h69D0] = 8'h06;
mem[16'h69D1] = 8'h6A;
mem[16'h69D2] = 8'h91;
mem[16'h69D3] = 8'h59;
mem[16'h69D4] = 8'hC8;
mem[16'h69D5] = 8'hA5;
mem[16'h69D6] = 8'h67;
mem[16'h69D7] = 8'h05;
mem[16'h69D8] = 8'h6D;
mem[16'h69D9] = 8'h51;
mem[16'h69DA] = 8'h59;
mem[16'h69DB] = 8'h5D;
mem[16'h69DC] = 8'h07;
mem[16'h69DD] = 8'h6A;
mem[16'h69DE] = 8'h91;
mem[16'h69DF] = 8'h59;
mem[16'h69E0] = 8'hC8;
mem[16'h69E1] = 8'hA5;
mem[16'h69E2] = 8'h68;
mem[16'h69E3] = 8'h05;
mem[16'h69E4] = 8'h6D;
mem[16'h69E5] = 8'h51;
mem[16'h69E6] = 8'h59;
mem[16'h69E7] = 8'h5D;
mem[16'h69E8] = 8'h08;
mem[16'h69E9] = 8'h6A;
mem[16'h69EA] = 8'h91;
mem[16'h69EB] = 8'h59;
mem[16'h69EC] = 8'hE6;
mem[16'h69ED] = 8'h56;
mem[16'h69EE] = 8'hA5;
mem[16'h69EF] = 8'h76;
mem[16'h69F0] = 8'h18;
mem[16'h69F1] = 8'h69;
mem[16'h69F2] = 8'h03;
mem[16'h69F3] = 8'h85;
mem[16'h69F4] = 8'h76;
mem[16'h69F5] = 8'hA6;
mem[16'h69F6] = 8'h62;
mem[16'h69F7] = 8'hE8;
mem[16'h69F8] = 8'hE0;
mem[16'h69F9] = 8'h1A;
mem[16'h69FA] = 8'hB0;
mem[16'h69FB] = 8'h03;
mem[16'h69FC] = 8'h4C;
mem[16'h69FD] = 8'h37;
mem[16'h69FE] = 8'h69;
mem[16'h69FF] = 8'hA5;
mem[16'h6A00] = 8'h77;
mem[16'h6A01] = 8'h49;
mem[16'h6A02] = 8'h01;
mem[16'h6A03] = 8'h85;
mem[16'h6A04] = 8'h77;
mem[16'h6A05] = 8'h60;
mem[16'h6A06] = 8'h2A;
mem[16'h6A07] = 8'h10;
mem[16'h6A08] = 8'h00;
mem[16'h6A09] = 8'h0A;
mem[16'h6A0A] = 8'h55;
mem[16'h6A0B] = 8'h00;
mem[16'h6A0C] = 8'h08;
mem[16'h6A0D] = 8'h54;
mem[16'h6A0E] = 8'h00;
mem[16'h6A0F] = 8'h2A;
mem[16'h6A10] = 8'h44;
mem[16'h6A11] = 8'h00;
mem[16'h6A12] = 8'h2A;
mem[16'h6A13] = 8'h51;
mem[16'h6A14] = 8'h00;
mem[16'h6A15] = 8'h0A;
mem[16'h6A16] = 8'h55;
mem[16'h6A17] = 8'h00;
mem[16'h6A18] = 8'h08;
mem[16'h6A19] = 8'h54;
mem[16'h6A1A] = 8'h00;
mem[16'h6A1B] = 8'h2A;
mem[16'h6A1C] = 8'h44;
mem[16'h6A1D] = 8'h00;
mem[16'h6A1E] = 8'h2A;
mem[16'h6A1F] = 8'h51;
mem[16'h6A20] = 8'h00;
mem[16'h6A21] = 8'h22;
mem[16'h6A22] = 8'h55;
mem[16'h6A23] = 8'h00;
mem[16'h6A24] = 8'h08;
mem[16'h6A25] = 8'h54;
mem[16'h6A26] = 8'h00;
mem[16'h6A27] = 8'h2A;
mem[16'h6A28] = 8'h44;
mem[16'h6A29] = 8'h00;
mem[16'h6A2A] = 8'h2A;
mem[16'h6A2B] = 8'h51;
mem[16'h6A2C] = 8'h00;
mem[16'h6A2D] = 8'h59;
mem[16'h6A2E] = 8'hE8;
mem[16'h6A2F] = 8'hE0;
mem[16'h6A30] = 8'hBE;
mem[16'h6A31] = 8'hD0;
mem[16'h6A32] = 8'hED;
mem[16'h6A33] = 8'h60;
mem[16'h6A34] = 8'hB1;
mem[16'h6A35] = 8'hAD;
mem[16'h6A36] = 8'hD0;
mem[16'h6A37] = 8'h4D;
mem[16'h6A38] = 8'hC9;
mem[16'h6A39] = 8'h4D;
mem[16'h6A3A] = 8'hD0;
mem[16'h6A3B] = 8'h44;
mem[16'h6A3C] = 8'hAE;
mem[16'h6A3D] = 8'hB0;
mem[16'h6A3E] = 8'h4A;
mem[16'h6A3F] = 8'hCA;
mem[16'h6A40] = 8'hE0;
mem[16'h6A41] = 8'h08;
mem[16'h6A42] = 8'h8D;
mem[16'h6A43] = 8'h59;
mem[16'h6A44] = 8'h69;
mem[16'h6A45] = 8'h8D;
mem[16'h6A46] = 8'h60;
mem[16'h6A47] = 8'h69;
mem[16'h6A48] = 8'h8D;
mem[16'h6A49] = 8'h68;
mem[16'h6A4A] = 8'h69;
mem[16'h6A4B] = 8'h8C;
mem[16'h6A4C] = 8'h5A;
mem[16'h6A4D] = 8'h69;
mem[16'h6A4E] = 8'h8C;
mem[16'h6A4F] = 8'h61;
mem[16'h6A50] = 8'h69;
mem[16'h6A51] = 8'h8C;
mem[16'h6A52] = 8'h69;
mem[16'h6A53] = 8'h69;
mem[16'h6A54] = 8'h60;
mem[16'h6A55] = 8'hA2;
mem[16'h6A56] = 8'h01;
mem[16'h6A57] = 8'h20;
mem[16'h6A58] = 8'h60;
mem[16'h6A59] = 8'h6A;
mem[16'h6A5A] = 8'hA2;
mem[16'h6A5B] = 8'h00;
mem[16'h6A5C] = 8'h20;
mem[16'h6A5D] = 8'h60;
mem[16'h6A5E] = 8'h6A;
mem[16'h6A5F] = 8'h60;
mem[16'h6A60] = 8'h86;
mem[16'h6A61] = 8'h70;
mem[16'h6A62] = 8'hBD;
mem[16'h6A63] = 8'hC2;
mem[16'h6A64] = 8'h62;
mem[16'h6A65] = 8'hD0;
mem[16'h6A66] = 8'h01;
mem[16'h6A67] = 8'h60;
mem[16'h6A68] = 8'hBD;
mem[16'h6A69] = 8'hBE;
mem[16'h6A6A] = 8'h62;
mem[16'h6A6B] = 8'hC9;
mem[16'h6A6C] = 8'h33;
mem[16'h6A6D] = 8'hF0;
mem[16'h6A6E] = 8'h23;
mem[16'h6A6F] = 8'hA5;
mem[16'h6A70] = 8'h8B;
mem[16'h6A71] = 8'hD0;
mem[16'h6A72] = 8'h10;
mem[16'h6A73] = 8'hBD;
mem[16'h6A74] = 8'hBC;
mem[16'h6A75] = 8'h62;
mem[16'h6A76] = 8'hC9;
mem[16'h6A77] = 8'h02;
mem[16'h6A78] = 8'h90;
mem[16'h6A79] = 8'h0A;
mem[16'h6A7A] = 8'h38;
mem[16'h6A7B] = 8'hE9;
mem[16'h6A7C] = 8'h02;
mem[16'h6A7D] = 8'h9D;
mem[16'h6A7E] = 8'hBC;
mem[16'h6A7F] = 8'h62;
mem[16'h6A80] = 8'h20;
mem[16'h6A81] = 8'h32;
mem[16'h6A82] = 8'h6C;
mem[16'h6A83] = 8'h60;
mem[16'h6A84] = 8'h20;
mem[16'h6A85] = 8'hC4;
mem[16'h6A86] = 8'h62;
mem[16'h6A87] = 8'hA9;
mem[16'h6A88] = 8'h00;
mem[16'h6A89] = 8'hA6;
mem[16'h6A8A] = 8'h70;
mem[16'h6A8B] = 8'h9D;
mem[16'h6A8C] = 8'hC2;
mem[16'h6A8D] = 8'h62;
mem[16'h6A8E] = 8'h8D;
mem[16'h6A8F] = 8'hD8;
mem[16'h6A90] = 8'h77;
mem[16'h6A91] = 8'h60;
mem[16'h6A92] = 8'hBD;
mem[16'h6A93] = 8'h07;
mem[16'h6A94] = 8'h6B;
mem[16'h6A95] = 8'h49;
mem[16'h6A96] = 8'h01;
mem[16'h6A97] = 8'h9D;
mem[16'h6A98] = 8'h07;
mem[16'h6A99] = 8'h6B;
mem[16'h6A9A] = 8'hF0;
mem[16'h6A9B] = 8'h4D;
mem[16'h6A9C] = 8'hBD;
mem[16'h6A9D] = 8'hBC;
mem[16'h6A9E] = 8'h62;
mem[16'h6A9F] = 8'h38;
mem[16'h6AA0] = 8'hED;
mem[16'h6AA1] = 8'h10;
mem[16'h6AA2] = 8'h51;
mem[16'h6AA3] = 8'h18;
mem[16'h6AA4] = 8'h6D;
mem[16'h6AA5] = 8'h16;
mem[16'h6AA6] = 8'h51;
mem[16'h6AA7] = 8'h20;
mem[16'h6AA8] = 8'h62;
mem[16'h6AA9] = 8'h65;
mem[16'h6AAA] = 8'hC9;
mem[16'h6AAB] = 8'h07;
mem[16'h6AAC] = 8'hB0;
mem[16'h6AAD] = 8'h3C;
mem[16'h6AAE] = 8'h20;
mem[16'h6AAF] = 8'hC4;
mem[16'h6AB0] = 8'h62;
mem[16'h6AB1] = 8'hA9;
mem[16'h6AB2] = 8'h00;
mem[16'h6AB3] = 8'hA6;
mem[16'h6AB4] = 8'h70;
mem[16'h6AB5] = 8'h9D;
mem[16'h6AB6] = 8'hC2;
mem[16'h6AB7] = 8'h62;
mem[16'h6AB8] = 8'h8D;
mem[16'h6AB9] = 8'hD9;
mem[16'h6ABA] = 8'h77;
mem[16'h6ABB] = 8'hA0;
mem[16'h6ABC] = 8'h00;
mem[16'h6ABD] = 8'hAD;
mem[16'h6ABE] = 8'hC0;
mem[16'h6ABF] = 8'h62;
mem[16'h6AC0] = 8'hF0;
mem[16'h6AC1] = 8'h07;
mem[16'h6AC2] = 8'hA0;
mem[16'h6AC3] = 8'h01;
mem[16'h6AC4] = 8'hAD;
mem[16'h6AC5] = 8'hC1;
mem[16'h6AC6] = 8'h62;
mem[16'h6AC7] = 8'hD0;
mem[16'h6AC8] = 8'h20;
mem[16'h6AC9] = 8'hAD;
mem[16'h6ACA] = 8'h13;
mem[16'h6ACB] = 8'h87;
mem[16'h6ACC] = 8'h29;
mem[16'h6ACD] = 8'h01;
mem[16'h6ACE] = 8'hF0;
mem[16'h6ACF] = 8'h19;
mem[16'h6AD0] = 8'hA9;
mem[16'h6AD1] = 8'h01;
mem[16'h6AD2] = 8'h8D;
mem[16'h6AD3] = 8'hD9;
mem[16'h6AD4] = 8'h77;
mem[16'h6AD5] = 8'h99;
mem[16'h6AD6] = 8'hC0;
mem[16'h6AD7] = 8'h62;
mem[16'h6AD8] = 8'hBD;
mem[16'h6AD9] = 8'hBE;
mem[16'h6ADA] = 8'h62;
mem[16'h6ADB] = 8'h99;
mem[16'h6ADC] = 8'hBA;
mem[16'h6ADD] = 8'h62;
mem[16'h6ADE] = 8'hBD;
mem[16'h6ADF] = 8'hBC;
mem[16'h6AE0] = 8'h62;
mem[16'h6AE1] = 8'h99;
mem[16'h6AE2] = 8'hB8;
mem[16'h6AE3] = 8'h62;
mem[16'h6AE4] = 8'h84;
mem[16'h6AE5] = 8'h70;
mem[16'h6AE6] = 8'h20;
mem[16'h6AE7] = 8'hF8;
mem[16'h6AE8] = 8'h62;
mem[16'h6AE9] = 8'h60;
mem[16'h6AEA] = 8'hBD;
mem[16'h6AEB] = 8'hBC;
mem[16'h6AEC] = 8'h62;
mem[16'h6AED] = 8'h38;
mem[16'h6AEE] = 8'hE9;
mem[16'h6AEF] = 8'h02;
mem[16'h6AF0] = 8'h90;
mem[16'h6AF1] = 8'h07;
mem[16'h6AF2] = 8'h9D;
mem[16'h6AF3] = 8'hBC;
mem[16'h6AF4] = 8'h62;
mem[16'h6AF5] = 8'h20;
mem[16'h6AF6] = 8'h32;
mem[16'h6AF7] = 8'h6C;
mem[16'h6AF8] = 8'h60;
mem[16'h6AF9] = 8'h20;
mem[16'h6AFA] = 8'hC4;
mem[16'h6AFB] = 8'h62;
mem[16'h6AFC] = 8'hA9;
mem[16'h6AFD] = 8'hEA;
mem[16'h6AFE] = 8'hA6;
mem[16'h6AFF] = 8'h70;
mem[16'h6B00] = 8'h9D;
mem[16'h6B01] = 8'hBC;
mem[16'h6B02] = 8'h62;
mem[16'h6B03] = 8'h20;
mem[16'h6B04] = 8'hC4;
mem[16'h6B05] = 8'h62;
mem[16'h6B06] = 8'h60;
mem[16'h6B07] = 8'h00;
mem[16'h6B08] = 8'h00;
mem[16'h6B09] = 8'hA2;
mem[16'h6B0A] = 8'h01;
mem[16'h6B0B] = 8'h20;
mem[16'h6B0C] = 8'h14;
mem[16'h6B0D] = 8'h6B;
mem[16'h6B0E] = 8'hA2;
mem[16'h6B0F] = 8'h00;
mem[16'h6B10] = 8'h20;
mem[16'h6B11] = 8'h14;
mem[16'h6B12] = 8'h6B;
mem[16'h6B13] = 8'h60;
mem[16'h6B14] = 8'h86;
mem[16'h6B15] = 8'h70;
mem[16'h6B16] = 8'hBD;
mem[16'h6B17] = 8'hC0;
mem[16'h6B18] = 8'h62;
mem[16'h6B19] = 8'hD0;
mem[16'h6B1A] = 8'h01;
mem[16'h6B1B] = 8'h60;
mem[16'h6B1C] = 8'hBD;
mem[16'h6B1D] = 8'hBA;
mem[16'h6B1E] = 8'h62;
mem[16'h6B1F] = 8'hC9;
mem[16'h6B20] = 8'h33;
mem[16'h6B21] = 8'hF0;
mem[16'h6B22] = 8'h24;
mem[16'h6B23] = 8'hA5;
mem[16'h6B24] = 8'h8B;
mem[16'h6B25] = 8'hD0;
mem[16'h6B26] = 8'h1F;
mem[16'h6B27] = 8'h20;
mem[16'h6B28] = 8'hFE;
mem[16'h6B29] = 8'h6B;
mem[16'h6B2A] = 8'hA6;
mem[16'h6B2B] = 8'h70;
mem[16'h6B2C] = 8'hBD;
mem[16'h6B2D] = 8'hB8;
mem[16'h6B2E] = 8'h62;
mem[16'h6B2F] = 8'h18;
mem[16'h6B30] = 8'h69;
mem[16'h6B31] = 8'h02;
mem[16'h6B32] = 8'h9D;
mem[16'h6B33] = 8'hB8;
mem[16'h6B34] = 8'h62;
mem[16'h6B35] = 8'hC9;
mem[16'h6B36] = 8'hEA;
mem[16'h6B37] = 8'h90;
mem[16'h6B38] = 8'h0D;
mem[16'h6B39] = 8'h20;
mem[16'h6B3A] = 8'hF8;
mem[16'h6B3B] = 8'h62;
mem[16'h6B3C] = 8'hA9;
mem[16'h6B3D] = 8'h00;
mem[16'h6B3E] = 8'hA6;
mem[16'h6B3F] = 8'h70;
mem[16'h6B40] = 8'h9D;
mem[16'h6B41] = 8'hC0;
mem[16'h6B42] = 8'h62;
mem[16'h6B43] = 8'h8D;
mem[16'h6B44] = 8'hD8;
mem[16'h6B45] = 8'h77;
mem[16'h6B46] = 8'h60;
mem[16'h6B47] = 8'hBD;
mem[16'h6B48] = 8'hB8;
mem[16'h6B49] = 8'h62;
mem[16'h6B4A] = 8'hC9;
mem[16'h6B4B] = 8'hEA;
mem[16'h6B4C] = 8'h90;
mem[16'h6B4D] = 8'h03;
mem[16'h6B4E] = 8'h4C;
mem[16'h6B4F] = 8'hEF;
mem[16'h6B50] = 8'h6B;
mem[16'h6B51] = 8'h20;
mem[16'h6B52] = 8'hFE;
mem[16'h6B53] = 8'h6B;
mem[16'h6B54] = 8'hA6;
mem[16'h6B55] = 8'h70;
mem[16'h6B56] = 8'hBD;
mem[16'h6B57] = 8'hB8;
mem[16'h6B58] = 8'h62;
mem[16'h6B59] = 8'h18;
mem[16'h6B5A] = 8'h69;
mem[16'h6B5B] = 8'h02;
mem[16'h6B5C] = 8'h9D;
mem[16'h6B5D] = 8'hB8;
mem[16'h6B5E] = 8'h62;
mem[16'h6B5F] = 8'h18;
mem[16'h6B60] = 8'h69;
mem[16'h6B61] = 8'h10;
mem[16'h6B62] = 8'h38;
mem[16'h6B63] = 8'hED;
mem[16'h6B64] = 8'h10;
mem[16'h6B65] = 8'h51;
mem[16'h6B66] = 8'h20;
mem[16'h6B67] = 8'h62;
mem[16'h6B68] = 8'h65;
mem[16'h6B69] = 8'hC9;
mem[16'h6B6A] = 8'h07;
mem[16'h6B6B] = 8'hB0;
mem[16'h6B6C] = 8'h38;
mem[16'h6B6D] = 8'h20;
mem[16'h6B6E] = 8'hF8;
mem[16'h6B6F] = 8'h62;
mem[16'h6B70] = 8'hA9;
mem[16'h6B71] = 8'h00;
mem[16'h6B72] = 8'hA6;
mem[16'h6B73] = 8'h70;
mem[16'h6B74] = 8'h9D;
mem[16'h6B75] = 8'hC0;
mem[16'h6B76] = 8'h62;
mem[16'h6B77] = 8'h8D;
mem[16'h6B78] = 8'hD9;
mem[16'h6B79] = 8'h77;
mem[16'h6B7A] = 8'hAC;
mem[16'h6B7B] = 8'hC7;
mem[16'h6B7C] = 8'h77;
mem[16'h6B7D] = 8'h88;
mem[16'h6B7E] = 8'hB9;
mem[16'h6B7F] = 8'hC2;
mem[16'h6B80] = 8'h62;
mem[16'h6B81] = 8'hD0;
mem[16'h6B82] = 8'h21;
mem[16'h6B83] = 8'hAD;
mem[16'h6B84] = 8'h14;
mem[16'h6B85] = 8'h87;
mem[16'h6B86] = 8'h6A;
mem[16'h6B87] = 8'h29;
mem[16'h6B88] = 8'h01;
mem[16'h6B89] = 8'hF0;
mem[16'h6B8A] = 8'h19;
mem[16'h6B8B] = 8'hA9;
mem[16'h6B8C] = 8'h01;
mem[16'h6B8D] = 8'h8D;
mem[16'h6B8E] = 8'hD9;
mem[16'h6B8F] = 8'h77;
mem[16'h6B90] = 8'h99;
mem[16'h6B91] = 8'hC2;
mem[16'h6B92] = 8'h62;
mem[16'h6B93] = 8'hBD;
mem[16'h6B94] = 8'hBA;
mem[16'h6B95] = 8'h62;
mem[16'h6B96] = 8'h99;
mem[16'h6B97] = 8'hBE;
mem[16'h6B98] = 8'h62;
mem[16'h6B99] = 8'hBD;
mem[16'h6B9A] = 8'hB8;
mem[16'h6B9B] = 8'h62;
mem[16'h6B9C] = 8'h99;
mem[16'h6B9D] = 8'hBC;
mem[16'h6B9E] = 8'h62;
mem[16'h6B9F] = 8'h84;
mem[16'h6BA0] = 8'h70;
mem[16'h6BA1] = 8'h20;
mem[16'h6BA2] = 8'hC4;
mem[16'h6BA3] = 8'h62;
mem[16'h6BA4] = 8'h60;
mem[16'h6BA5] = 8'hBD;
mem[16'h6BA6] = 8'hB8;
mem[16'h6BA7] = 8'h62;
mem[16'h6BA8] = 8'hC9;
mem[16'h6BA9] = 8'hEA;
mem[16'h6BAA] = 8'hB0;
mem[16'h6BAB] = 8'h43;
mem[16'h6BAC] = 8'h20;
mem[16'h6BAD] = 8'hFE;
mem[16'h6BAE] = 8'h6B;
mem[16'h6BAF] = 8'hA6;
mem[16'h6BB0] = 8'h70;
mem[16'h6BB1] = 8'hBD;
mem[16'h6BB2] = 8'hB8;
mem[16'h6BB3] = 8'h62;
mem[16'h6BB4] = 8'h18;
mem[16'h6BB5] = 8'h69;
mem[16'h6BB6] = 8'h02;
mem[16'h6BB7] = 8'h9D;
mem[16'h6BB8] = 8'hB8;
mem[16'h6BB9] = 8'h62;
mem[16'h6BBA] = 8'h18;
mem[16'h6BBB] = 8'h69;
mem[16'h6BBC] = 8'h10;
mem[16'h6BBD] = 8'h38;
mem[16'h6BBE] = 8'hED;
mem[16'h6BBF] = 8'h10;
mem[16'h6BC0] = 8'h51;
mem[16'h6BC1] = 8'h20;
mem[16'h6BC2] = 8'h62;
mem[16'h6BC3] = 8'h65;
mem[16'h6BC4] = 8'hC9;
mem[16'h6BC5] = 8'h07;
mem[16'h6BC6] = 8'h90;
mem[16'h6BC7] = 8'hA5;
mem[16'h6BC8] = 8'hBD;
mem[16'h6BC9] = 8'hB8;
mem[16'h6BCA] = 8'h62;
mem[16'h6BCB] = 8'hC9;
mem[16'h6BCC] = 8'hEA;
mem[16'h6BCD] = 8'hB0;
mem[16'h6BCE] = 8'h20;
mem[16'h6BCF] = 8'h20;
mem[16'h6BD0] = 8'hFE;
mem[16'h6BD1] = 8'h6B;
mem[16'h6BD2] = 8'hA6;
mem[16'h6BD3] = 8'h70;
mem[16'h6BD4] = 8'hBD;
mem[16'h6BD5] = 8'hB8;
mem[16'h6BD6] = 8'h62;
mem[16'h6BD7] = 8'h18;
mem[16'h6BD8] = 8'h69;
mem[16'h6BD9] = 8'h02;
mem[16'h6BDA] = 8'h9D;
mem[16'h6BDB] = 8'hB8;
mem[16'h6BDC] = 8'h62;
mem[16'h6BDD] = 8'h18;
mem[16'h6BDE] = 8'h69;
mem[16'h6BDF] = 8'h10;
mem[16'h6BE0] = 8'h38;
mem[16'h6BE1] = 8'hED;
mem[16'h6BE2] = 8'h10;
mem[16'h6BE3] = 8'h51;
mem[16'h6BE4] = 8'h20;
mem[16'h6BE5] = 8'h62;
mem[16'h6BE6] = 8'h65;
mem[16'h6BE7] = 8'hC9;
mem[16'h6BE8] = 8'h07;
mem[16'h6BE9] = 8'hB0;
mem[16'h6BEA] = 8'h03;
mem[16'h6BEB] = 8'h4C;
mem[16'h6BEC] = 8'h6D;
mem[16'h6BED] = 8'h6B;
mem[16'h6BEE] = 8'h60;
mem[16'h6BEF] = 8'h20;
mem[16'h6BF0] = 8'hF8;
mem[16'h6BF1] = 8'h62;
mem[16'h6BF2] = 8'hA9;
mem[16'h6BF3] = 8'h01;
mem[16'h6BF4] = 8'hA6;
mem[16'h6BF5] = 8'h70;
mem[16'h6BF6] = 8'h9D;
mem[16'h6BF7] = 8'hB8;
mem[16'h6BF8] = 8'h62;
mem[16'h6BF9] = 8'h20;
mem[16'h6BFA] = 8'hF8;
mem[16'h6BFB] = 8'h62;
mem[16'h6BFC] = 8'h60;
mem[16'h6BFD] = 8'h00;
mem[16'h6BFE] = 8'hA6;
mem[16'h6BFF] = 8'h70;
mem[16'h6C00] = 8'hBD;
mem[16'h6C01] = 8'hBA;
mem[16'h6C02] = 8'h62;
mem[16'h6C03] = 8'h85;
mem[16'h6C04] = 8'h56;
mem[16'h6C05] = 8'hBC;
mem[16'h6C06] = 8'hB8;
mem[16'h6C07] = 8'h62;
mem[16'h6C08] = 8'h84;
mem[16'h6C09] = 8'h57;
mem[16'h6C0A] = 8'hB9;
mem[16'h6C0B] = 8'h3E;
mem[16'h6C0C] = 8'h8C;
mem[16'h6C0D] = 8'hAA;
mem[16'h6C0E] = 8'hBD;
mem[16'h6C0F] = 8'h94;
mem[16'h6C10] = 8'h8E;
mem[16'h6C11] = 8'hAA;
mem[16'h6C12] = 8'hBD;
mem[16'h6C13] = 8'h24;
mem[16'h6C14] = 8'h6C;
mem[16'h6C15] = 8'hBC;
mem[16'h6C16] = 8'h2B;
mem[16'h6C17] = 8'h6C;
mem[16'h6C18] = 8'h20;
mem[16'h6C19] = 8'hD1;
mem[16'h6C1A] = 8'h8A;
mem[16'h6C1B] = 8'hA9;
mem[16'h6C1C] = 8'h20;
mem[16'h6C1D] = 8'h8D;
mem[16'h6C1E] = 8'hCA;
mem[16'h6C1F] = 8'h8A;
mem[16'h6C20] = 8'h20;
mem[16'h6C21] = 8'h79;
mem[16'h6C22] = 8'h8A;
mem[16'h6C23] = 8'h60;
mem[16'h6C24] = 8'h66;
mem[16'h6C25] = 8'h86;
mem[16'h6C26] = 8'hA6;
mem[16'h6C27] = 8'hC6;
mem[16'h6C28] = 8'hE6;
mem[16'h6C29] = 8'h06;
mem[16'h6C2A] = 8'h26;
mem[16'h6C2B] = 8'h6C;
mem[16'h6C2C] = 8'h6C;
mem[16'h6C2D] = 8'h6C;
mem[16'h6C2E] = 8'h6C;
mem[16'h6C2F] = 8'h6C;
mem[16'h6C30] = 8'h6D;
mem[16'h6C31] = 8'h6D;
mem[16'h6C32] = 8'hA6;
mem[16'h6C33] = 8'h70;
mem[16'h6C34] = 8'hBD;
mem[16'h6C35] = 8'hBE;
mem[16'h6C36] = 8'h62;
mem[16'h6C37] = 8'h85;
mem[16'h6C38] = 8'h56;
mem[16'h6C39] = 8'hBC;
mem[16'h6C3A] = 8'hBC;
mem[16'h6C3B] = 8'h62;
mem[16'h6C3C] = 8'h84;
mem[16'h6C3D] = 8'h57;
mem[16'h6C3E] = 8'hB9;
mem[16'h6C3F] = 8'h3E;
mem[16'h6C40] = 8'h8C;
mem[16'h6C41] = 8'hAA;
mem[16'h6C42] = 8'hBD;
mem[16'h6C43] = 8'h94;
mem[16'h6C44] = 8'h8E;
mem[16'h6C45] = 8'hAA;
mem[16'h6C46] = 8'hBD;
mem[16'h6C47] = 8'h58;
mem[16'h6C48] = 8'h6C;
mem[16'h6C49] = 8'hBC;
mem[16'h6C4A] = 8'h5F;
mem[16'h6C4B] = 8'h6C;
mem[16'h6C4C] = 8'h20;
mem[16'h6C4D] = 8'hD1;
mem[16'h6C4E] = 8'h8A;
mem[16'h6C4F] = 8'hA9;
mem[16'h6C50] = 8'h20;
mem[16'h6C51] = 8'h8D;
mem[16'h6C52] = 8'hCA;
mem[16'h6C53] = 8'h8A;
mem[16'h6C54] = 8'h20;
mem[16'h6C55] = 8'h79;
mem[16'h6C56] = 8'h8A;
mem[16'h6C57] = 8'h60;
mem[16'h6C58] = 8'h93;
mem[16'h6C59] = 8'hB3;
mem[16'h6C5A] = 8'hD3;
mem[16'h6C5B] = 8'hF3;
mem[16'h6C5C] = 8'h13;
mem[16'h6C5D] = 8'h33;
mem[16'h6C5E] = 8'h53;
mem[16'h6C5F] = 8'h74;
mem[16'h6C60] = 8'h74;
mem[16'h6C61] = 8'h74;
mem[16'h6C62] = 8'h74;
mem[16'h6C63] = 8'h75;
mem[16'h6C64] = 8'h75;
mem[16'h6C65] = 8'h75;
mem[16'h6C66] = 8'h00;
mem[16'h6C67] = 8'h40;
mem[16'h6C68] = 8'h5D;
mem[16'h6C69] = 8'h00;
mem[16'h6C6A] = 8'h00;
mem[16'h6C6B] = 8'h60;
mem[16'h6C6C] = 8'h35;
mem[16'h6C6D] = 8'h00;
mem[16'h6C6E] = 8'h00;
mem[16'h6C6F] = 8'h60;
mem[16'h6C70] = 8'h06;
mem[16'h6C71] = 8'h00;
mem[16'h6C72] = 8'h78;
mem[16'h6C73] = 8'h60;
mem[16'h6C74] = 8'h03;
mem[16'h6C75] = 8'h00;
mem[16'h6C76] = 8'h4C;
mem[16'h6C77] = 8'h71;
mem[16'h6C78] = 8'h01;
mem[16'h6C79] = 8'h00;
mem[16'h6C7A] = 8'h7E;
mem[16'h6C7B] = 8'h7B;
mem[16'h6C7C] = 8'h00;
mem[16'h6C7D] = 8'h00;
mem[16'h6C7E] = 8'h4F;
mem[16'h6C7F] = 8'h31;
mem[16'h6C80] = 8'h00;
mem[16'h6C81] = 8'h00;
mem[16'h6C82] = 8'h05;
mem[16'h6C83] = 8'h1B;
mem[16'h6C84] = 8'h00;
mem[16'h6C85] = 8'h00;
mem[16'h6C86] = 8'h00;
mem[16'h6C87] = 8'h00;
mem[16'h6C88] = 8'h3B;
mem[16'h6C89] = 8'h01;
mem[16'h6C8A] = 8'h00;
mem[16'h6C8B] = 8'h40;
mem[16'h6C8C] = 8'h6B;
mem[16'h6C8D] = 8'h00;
mem[16'h6C8E] = 8'h00;
mem[16'h6C8F] = 8'h40;
mem[16'h6C90] = 8'h0D;
mem[16'h6C91] = 8'h00;
mem[16'h6C92] = 8'h70;
mem[16'h6C93] = 8'h41;
mem[16'h6C94] = 8'h07;
mem[16'h6C95] = 8'h00;
mem[16'h6C96] = 8'h18;
mem[16'h6C97] = 8'h63;
mem[16'h6C98] = 8'h03;
mem[16'h6C99] = 8'h00;
mem[16'h6C9A] = 8'h7C;
mem[16'h6C9B] = 8'h77;
mem[16'h6C9C] = 8'h01;
mem[16'h6C9D] = 8'h00;
mem[16'h6C9E] = 8'h1E;
mem[16'h6C9F] = 8'h63;
mem[16'h6CA0] = 8'h00;
mem[16'h6CA1] = 8'h00;
mem[16'h6CA2] = 8'h0A;
mem[16'h6CA3] = 8'h36;
mem[16'h6CA4] = 8'h00;
mem[16'h6CA5] = 8'h00;
mem[16'h6CA6] = 8'h00;
mem[16'h6CA7] = 8'h00;
mem[16'h6CA8] = 8'h76;
mem[16'h6CA9] = 8'h02;
mem[16'h6CAA] = 8'h00;
mem[16'h6CAB] = 8'h00;
mem[16'h6CAC] = 8'h57;
mem[16'h6CAD] = 8'h01;
mem[16'h6CAE] = 8'h00;
mem[16'h6CAF] = 8'h00;
mem[16'h6CB0] = 8'h1B;
mem[16'h6CB1] = 8'h00;
mem[16'h6CB2] = 8'h60;
mem[16'h6CB3] = 8'h03;
mem[16'h6CB4] = 8'h0F;
mem[16'h6CB5] = 8'h00;
mem[16'h6CB6] = 8'h30;
mem[16'h6CB7] = 8'h46;
mem[16'h6CB8] = 8'h07;
mem[16'h6CB9] = 8'h00;
mem[16'h6CBA] = 8'h78;
mem[16'h6CBB] = 8'h6F;
mem[16'h6CBC] = 8'h03;
mem[16'h6CBD] = 8'h00;
mem[16'h6CBE] = 8'h3C;
mem[16'h6CBF] = 8'h46;
mem[16'h6CC0] = 8'h01;
mem[16'h6CC1] = 8'h00;
mem[16'h6CC2] = 8'h14;
mem[16'h6CC3] = 8'h6C;
mem[16'h6CC4] = 8'h00;
mem[16'h6CC5] = 8'h00;
mem[16'h6CC6] = 8'h00;
mem[16'h6CC7] = 8'h00;
mem[16'h6CC8] = 8'h6C;
mem[16'h6CC9] = 8'h05;
mem[16'h6CCA] = 8'h00;
mem[16'h6CCB] = 8'h00;
mem[16'h6CCC] = 8'h2E;
mem[16'h6CCD] = 8'h03;
mem[16'h6CCE] = 8'h00;
mem[16'h6CCF] = 8'h00;
mem[16'h6CD0] = 8'h36;
mem[16'h6CD1] = 8'h00;
mem[16'h6CD2] = 8'h40;
mem[16'h6CD3] = 8'h07;
mem[16'h6CD4] = 8'h1E;
mem[16'h6CD5] = 8'h00;
mem[16'h6CD6] = 8'h60;
mem[16'h6CD7] = 8'h0C;
mem[16'h6CD8] = 8'h0F;
mem[16'h6CD9] = 8'h00;
mem[16'h6CDA] = 8'h70;
mem[16'h6CDB] = 8'h5F;
mem[16'h6CDC] = 8'h07;
mem[16'h6CDD] = 8'h00;
mem[16'h6CDE] = 8'h78;
mem[16'h6CDF] = 8'h0C;
mem[16'h6CE0] = 8'h03;
mem[16'h6CE1] = 8'h00;
mem[16'h6CE2] = 8'h28;
mem[16'h6CE3] = 8'h58;
mem[16'h6CE4] = 8'h01;
mem[16'h6CE5] = 8'h00;
mem[16'h6CE6] = 8'h00;
mem[16'h6CE7] = 8'h00;
mem[16'h6CE8] = 8'h58;
mem[16'h6CE9] = 8'h0B;
mem[16'h6CEA] = 8'h00;
mem[16'h6CEB] = 8'h00;
mem[16'h6CEC] = 8'h5C;
mem[16'h6CED] = 8'h06;
mem[16'h6CEE] = 8'h00;
mem[16'h6CEF] = 8'h00;
mem[16'h6CF0] = 8'h6C;
mem[16'h6CF1] = 8'h00;
mem[16'h6CF2] = 8'h00;
mem[16'h6CF3] = 8'h0F;
mem[16'h6CF4] = 8'h3C;
mem[16'h6CF5] = 8'h00;
mem[16'h6CF6] = 8'h40;
mem[16'h6CF7] = 8'h19;
mem[16'h6CF8] = 8'h1E;
mem[16'h6CF9] = 8'h00;
mem[16'h6CFA] = 8'h60;
mem[16'h6CFB] = 8'h3F;
mem[16'h6CFC] = 8'h0F;
mem[16'h6CFD] = 8'h00;
mem[16'h6CFE] = 8'h70;
mem[16'h6CFF] = 8'h19;
mem[16'h6D00] = 8'h06;
mem[16'h6D01] = 8'h00;
mem[16'h6D02] = 8'h50;
mem[16'h6D03] = 8'h30;
mem[16'h6D04] = 8'h03;
mem[16'h6D05] = 8'h00;
mem[16'h6D06] = 8'h00;
mem[16'h6D07] = 8'h00;
mem[16'h6D08] = 8'h30;
mem[16'h6D09] = 8'h17;
mem[16'h6D0A] = 8'h00;
mem[16'h6D0B] = 8'h00;
mem[16'h6D0C] = 8'h38;
mem[16'h6D0D] = 8'h0D;
mem[16'h6D0E] = 8'h00;
mem[16'h6D0F] = 8'h00;
mem[16'h6D10] = 8'h58;
mem[16'h6D11] = 8'h01;
mem[16'h6D12] = 8'h00;
mem[16'h6D13] = 8'h1E;
mem[16'h6D14] = 8'h78;
mem[16'h6D15] = 8'h00;
mem[16'h6D16] = 8'h00;
mem[16'h6D17] = 8'h33;
mem[16'h6D18] = 8'h3C;
mem[16'h6D19] = 8'h00;
mem[16'h6D1A] = 8'h40;
mem[16'h6D1B] = 8'h7F;
mem[16'h6D1C] = 8'h1E;
mem[16'h6D1D] = 8'h00;
mem[16'h6D1E] = 8'h60;
mem[16'h6D1F] = 8'h33;
mem[16'h6D20] = 8'h0C;
mem[16'h6D21] = 8'h00;
mem[16'h6D22] = 8'h20;
mem[16'h6D23] = 8'h61;
mem[16'h6D24] = 8'h06;
mem[16'h6D25] = 8'h00;
mem[16'h6D26] = 8'h00;
mem[16'h6D27] = 8'h00;
mem[16'h6D28] = 8'h60;
mem[16'h6D29] = 8'h2E;
mem[16'h6D2A] = 8'h00;
mem[16'h6D2B] = 8'h00;
mem[16'h6D2C] = 8'h70;
mem[16'h6D2D] = 8'h1A;
mem[16'h6D2E] = 8'h00;
mem[16'h6D2F] = 8'h00;
mem[16'h6D30] = 8'h30;
mem[16'h6D31] = 8'h03;
mem[16'h6D32] = 8'h00;
mem[16'h6D33] = 8'h3C;
mem[16'h6D34] = 8'h70;
mem[16'h6D35] = 8'h01;
mem[16'h6D36] = 8'h00;
mem[16'h6D37] = 8'h66;
mem[16'h6D38] = 8'h78;
mem[16'h6D39] = 8'h00;
mem[16'h6D3A] = 8'h00;
mem[16'h6D3B] = 8'h7F;
mem[16'h6D3C] = 8'h3D;
mem[16'h6D3D] = 8'h00;
mem[16'h6D3E] = 8'h40;
mem[16'h6D3F] = 8'h67;
mem[16'h6D40] = 8'h18;
mem[16'h6D41] = 8'h00;
mem[16'h6D42] = 8'h40;
mem[16'h6D43] = 8'h42;
mem[16'h6D44] = 8'h0D;
mem[16'h6D45] = 8'h00;
mem[16'h6D46] = 8'h20;
mem[16'h6D47] = 8'hBE;
mem[16'h6D48] = 8'h7E;
mem[16'h6D49] = 8'hAD;
mem[16'h6D4A] = 8'hC0;
mem[16'h6D4B] = 8'h62;
mem[16'h6D4C] = 8'hF0;
mem[16'h6D4D] = 8'h07;
mem[16'h6D4E] = 8'hA9;
mem[16'h6D4F] = 8'h00;
mem[16'h6D50] = 8'h85;
mem[16'h6D51] = 8'h70;
mem[16'h6D52] = 8'h20;
mem[16'h6D53] = 8'hF8;
mem[16'h6D54] = 8'h62;
mem[16'h6D55] = 8'hAD;
mem[16'h6D56] = 8'hC2;
mem[16'h6D57] = 8'h62;
mem[16'h6D58] = 8'hF0;
mem[16'h6D59] = 8'h07;
mem[16'h6D5A] = 8'hA9;
mem[16'h6D5B] = 8'h00;
mem[16'h6D5C] = 8'h85;
mem[16'h6D5D] = 8'h70;
mem[16'h6D5E] = 8'h20;
mem[16'h6D5F] = 8'hC4;
mem[16'h6D60] = 8'h62;
mem[16'h6D61] = 8'hA9;
mem[16'h6D62] = 8'h0A;
mem[16'h6D63] = 8'h8D;
mem[16'h6D64] = 8'hA5;
mem[16'h6D65] = 8'h71;
mem[16'h6D66] = 8'hA9;
mem[16'h6D67] = 8'h5B;
mem[16'h6D68] = 8'h85;
mem[16'h6D69] = 8'h57;
mem[16'h6D6A] = 8'hA9;
mem[16'h6D6B] = 8'h5E;
mem[16'h6D6C] = 8'h85;
mem[16'h6D6D] = 8'h56;
mem[16'h6D6E] = 8'h20;
mem[16'h6D6F] = 8'h5E;
mem[16'h6D70] = 8'h71;
mem[16'h6D71] = 8'hA5;
mem[16'h6D72] = 8'h57;
mem[16'h6D73] = 8'h18;
mem[16'h6D74] = 8'h69;
mem[16'h6D75] = 8'h08;
mem[16'h6D76] = 8'h85;
mem[16'h6D77] = 8'h57;
mem[16'h6D78] = 8'hC9;
mem[16'h6D79] = 8'hAF;
mem[16'h6D7A] = 8'h90;
mem[16'h6D7B] = 8'hEE;
mem[16'h6D7C] = 8'hA9;
mem[16'h6D7D] = 8'h0C;
mem[16'h6D7E] = 8'h85;
mem[16'h6D7F] = 8'h25;
mem[16'h6D80] = 8'hA9;
mem[16'h6D81] = 8'h0E;
mem[16'h6D82] = 8'h85;
mem[16'h6D83] = 8'h24;
mem[16'h6D84] = 8'hA9;
mem[16'h6D85] = 8'h9A;
mem[16'h6D86] = 8'h85;
mem[16'h6D87] = 8'h59;
mem[16'h6D88] = 8'hA9;
mem[16'h6D89] = 8'h6D;
mem[16'h6D8A] = 8'h85;
mem[16'h6D8B] = 8'h5A;
mem[16'h6D8C] = 8'h20;
mem[16'h6D8D] = 8'hD5;
mem[16'h6D8E] = 8'h67;
mem[16'h6D8F] = 8'h60;
mem[16'h6D90] = 8'h55;
mem[16'h6D91] = 8'h55;
mem[16'h6D92] = 8'h55;
mem[16'h6D93] = 8'h55;
mem[16'h6D94] = 8'h55;
mem[16'h6D95] = 8'h55;
mem[16'h6D96] = 8'h55;
mem[16'h6D97] = 8'h55;
mem[16'h6D98] = 8'h55;
mem[16'h6D99] = 8'h55;
mem[16'h6D9A] = 8'hA0;
mem[16'h6D9B] = 8'hC7;
mem[16'h6D9C] = 8'hC1;
mem[16'h6D9D] = 8'hCD;
mem[16'h6D9E] = 8'hC5;
mem[16'h6D9F] = 8'hA0;
mem[16'h6DA0] = 8'hCF;
mem[16'h6DA1] = 8'hD6;
mem[16'h6DA2] = 8'hC5;
mem[16'h6DA3] = 8'hD2;
mem[16'h6DA4] = 8'hA0;
mem[16'h6DA5] = 8'h00;
mem[16'h6DA6] = 8'hAD;
mem[16'h6DA7] = 8'hC0;
mem[16'h6DA8] = 8'h62;
mem[16'h6DA9] = 8'hF0;
mem[16'h6DAA] = 8'h07;
mem[16'h6DAB] = 8'hA9;
mem[16'h6DAC] = 8'h00;
mem[16'h6DAD] = 8'h85;
mem[16'h6DAE] = 8'h70;
mem[16'h6DAF] = 8'h20;
mem[16'h6DB0] = 8'hF8;
mem[16'h6DB1] = 8'h62;
mem[16'h6DB2] = 8'hAD;
mem[16'h6DB3] = 8'hC2;
mem[16'h6DB4] = 8'h62;
mem[16'h6DB5] = 8'hF0;
mem[16'h6DB6] = 8'h07;
mem[16'h6DB7] = 8'hA9;
mem[16'h6DB8] = 8'h00;
mem[16'h6DB9] = 8'h85;
mem[16'h6DBA] = 8'h70;
mem[16'h6DBB] = 8'h20;
mem[16'h6DBC] = 8'hC4;
mem[16'h6DBD] = 8'h62;
mem[16'h6DBE] = 8'hA9;
mem[16'h6DBF] = 8'h0A;
mem[16'h6DC0] = 8'h8D;
mem[16'h6DC1] = 8'hA5;
mem[16'h6DC2] = 8'h71;
mem[16'h6DC3] = 8'hA9;
mem[16'h6DC4] = 8'h5B;
mem[16'h6DC5] = 8'h85;
mem[16'h6DC6] = 8'h57;
mem[16'h6DC7] = 8'hA9;
mem[16'h6DC8] = 8'h5E;
mem[16'h6DC9] = 8'h85;
mem[16'h6DCA] = 8'h56;
mem[16'h6DCB] = 8'h20;
mem[16'h6DCC] = 8'h5E;
mem[16'h6DCD] = 8'h71;
mem[16'h6DCE] = 8'hA5;
mem[16'h6DCF] = 8'h57;
mem[16'h6DD0] = 8'h18;
mem[16'h6DD1] = 8'h69;
mem[16'h6DD2] = 8'h08;
mem[16'h6DD3] = 8'h85;
mem[16'h6DD4] = 8'h57;
mem[16'h6DD5] = 8'hC9;
mem[16'h6DD6] = 8'hB0;
mem[16'h6DD7] = 8'h90;
mem[16'h6DD8] = 8'hEE;
mem[16'h6DD9] = 8'hA9;
mem[16'h6DDA] = 8'h0C;
mem[16'h6DDB] = 8'h85;
mem[16'h6DDC] = 8'h25;
mem[16'h6DDD] = 8'hA9;
mem[16'h6DDE] = 8'h0E;
mem[16'h6DDF] = 8'h85;
mem[16'h6DE0] = 8'h24;
mem[16'h6DE1] = 8'hA9;
mem[16'h6DE2] = 8'h37;
mem[16'h6DE3] = 8'h85;
mem[16'h6DE4] = 8'h59;
mem[16'h6DE5] = 8'hA9;
mem[16'h6DE6] = 8'h6E;
mem[16'h6DE7] = 8'h85;
mem[16'h6DE8] = 8'h5A;
mem[16'h6DE9] = 8'h20;
mem[16'h6DEA] = 8'hD5;
mem[16'h6DEB] = 8'h67;
mem[16'h6DEC] = 8'h60;
mem[16'h6DED] = 8'hA9;
mem[16'h6DEE] = 8'h0C;
mem[16'h6DEF] = 8'h85;
mem[16'h6DF0] = 8'h25;
mem[16'h6DF1] = 8'hA9;
mem[16'h6DF2] = 8'h0E;
mem[16'h6DF3] = 8'h85;
mem[16'h6DF4] = 8'h24;
mem[16'h6DF5] = 8'hA9;
mem[16'h6DF6] = 8'h37;
mem[16'h6DF7] = 8'h85;
mem[16'h6DF8] = 8'h59;
mem[16'h6DF9] = 8'hA9;
mem[16'h6DFA] = 8'h6E;
mem[16'h6DFB] = 8'h85;
mem[16'h6DFC] = 8'h5A;
mem[16'h6DFD] = 8'h20;
mem[16'h6DFE] = 8'hD5;
mem[16'h6DFF] = 8'h67;
mem[16'h6E00] = 8'hA9;
mem[16'h6E01] = 8'h5B;
mem[16'h6E02] = 8'h8D;
mem[16'h6E03] = 8'hA1;
mem[16'h6E04] = 8'h55;
mem[16'h6E05] = 8'hA9;
mem[16'h6E06] = 8'h5E;
mem[16'h6E07] = 8'h8D;
mem[16'h6E08] = 8'hA2;
mem[16'h6E09] = 8'h55;
mem[16'h6E0A] = 8'h20;
mem[16'h6E0B] = 8'h51;
mem[16'h6E0C] = 8'h55;
mem[16'h6E0D] = 8'hA9;
mem[16'h6E0E] = 8'h63;
mem[16'h6E0F] = 8'h8D;
mem[16'h6E10] = 8'hA2;
mem[16'h6E11] = 8'h55;
mem[16'h6E12] = 8'h20;
mem[16'h6E13] = 8'h51;
mem[16'h6E14] = 8'h55;
mem[16'h6E15] = 8'hAD;
mem[16'h6E16] = 8'hA1;
mem[16'h6E17] = 8'h55;
mem[16'h6E18] = 8'h18;
mem[16'h6E19] = 8'h69;
mem[16'h6E1A] = 8'h08;
mem[16'h6E1B] = 8'h8D;
mem[16'h6E1C] = 8'hA1;
mem[16'h6E1D] = 8'h55;
mem[16'h6E1E] = 8'hC9;
mem[16'h6E1F] = 8'hB0;
mem[16'h6E20] = 8'h90;
mem[16'h6E21] = 8'hE3;
mem[16'h6E22] = 8'hA9;
mem[16'h6E23] = 8'h00;
mem[16'h6E24] = 8'h85;
mem[16'h6E25] = 8'h70;
mem[16'h6E26] = 8'hAD;
mem[16'h6E27] = 8'hC0;
mem[16'h6E28] = 8'h62;
mem[16'h6E29] = 8'hF0;
mem[16'h6E2A] = 8'h03;
mem[16'h6E2B] = 8'h20;
mem[16'h6E2C] = 8'hF8;
mem[16'h6E2D] = 8'h62;
mem[16'h6E2E] = 8'hAD;
mem[16'h6E2F] = 8'hC2;
mem[16'h6E30] = 8'h62;
mem[16'h6E31] = 8'hF0;
mem[16'h6E32] = 8'h03;
mem[16'h6E33] = 8'h20;
mem[16'h6E34] = 8'hC4;
mem[16'h6E35] = 8'h62;
mem[16'h6E36] = 8'h60;
mem[16'h6E37] = 8'hA0;
mem[16'h6E38] = 8'hD4;
mem[16'h6E39] = 8'hC9;
mem[16'h6E3A] = 8'hCD;
mem[16'h6E3B] = 8'hC5;
mem[16'h6E3C] = 8'hA0;
mem[16'h6E3D] = 8'hCF;
mem[16'h6E3E] = 8'hD6;
mem[16'h6E3F] = 8'hC5;
mem[16'h6E40] = 8'hD2;
mem[16'h6E41] = 8'hA0;
mem[16'h6E42] = 8'h00;
mem[16'h6E43] = 8'hAD;
mem[16'h6E44] = 8'hC0;
mem[16'h6E45] = 8'h62;
mem[16'h6E46] = 8'hF0;
mem[16'h6E47] = 8'h07;
mem[16'h6E48] = 8'hA9;
mem[16'h6E49] = 8'h00;
mem[16'h6E4A] = 8'h85;
mem[16'h6E4B] = 8'h70;
mem[16'h6E4C] = 8'h20;
mem[16'h6E4D] = 8'hF8;
mem[16'h6E4E] = 8'h62;
mem[16'h6E4F] = 8'hAD;
mem[16'h6E50] = 8'hC2;
mem[16'h6E51] = 8'h62;
mem[16'h6E52] = 8'hF0;
mem[16'h6E53] = 8'h07;
mem[16'h6E54] = 8'hA2;
mem[16'h6E55] = 8'h00;
mem[16'h6E56] = 8'h86;
mem[16'h6E57] = 8'h70;
mem[16'h6E58] = 8'h20;
mem[16'h6E59] = 8'hC4;
mem[16'h6E5A] = 8'h62;
mem[16'h6E5B] = 8'hA9;
mem[16'h6E5C] = 8'h0A;
mem[16'h6E5D] = 8'h8D;
mem[16'h6E5E] = 8'hA5;
mem[16'h6E5F] = 8'h71;
mem[16'h6E60] = 8'hA9;
mem[16'h6E61] = 8'h61;
mem[16'h6E62] = 8'h85;
mem[16'h6E63] = 8'h57;
mem[16'h6E64] = 8'hA9;
mem[16'h6E65] = 8'h5E;
mem[16'h6E66] = 8'h85;
mem[16'h6E67] = 8'h56;
mem[16'h6E68] = 8'h20;
mem[16'h6E69] = 8'h5E;
mem[16'h6E6A] = 8'h71;
mem[16'h6E6B] = 8'hA5;
mem[16'h6E6C] = 8'h57;
mem[16'h6E6D] = 8'h18;
mem[16'h6E6E] = 8'h69;
mem[16'h6E6F] = 8'h08;
mem[16'h6E70] = 8'h85;
mem[16'h6E71] = 8'h57;
mem[16'h6E72] = 8'hC9;
mem[16'h6E73] = 8'hA8;
mem[16'h6E74] = 8'h90;
mem[16'h6E75] = 8'hEE;
mem[16'h6E76] = 8'hA9;
mem[16'h6E77] = 8'h0C;
mem[16'h6E78] = 8'h85;
mem[16'h6E79] = 8'h25;
mem[16'h6E7A] = 8'hA9;
mem[16'h6E7B] = 8'h0F;
mem[16'h6E7C] = 8'h85;
mem[16'h6E7D] = 8'h24;
mem[16'h6E7E] = 8'hA9;
mem[16'h6E7F] = 8'hF1;
mem[16'h6E80] = 8'h85;
mem[16'h6E81] = 8'h59;
mem[16'h6E82] = 8'hA9;
mem[16'h6E83] = 8'h6E;
mem[16'h6E84] = 8'h85;
mem[16'h6E85] = 8'h5A;
mem[16'h6E86] = 8'h20;
mem[16'h6E87] = 8'hD5;
mem[16'h6E88] = 8'h67;
mem[16'h6E89] = 8'hA9;
mem[16'h6E8A] = 8'h0C;
mem[16'h6E8B] = 8'h85;
mem[16'h6E8C] = 8'h25;
mem[16'h6E8D] = 8'hA9;
mem[16'h6E8E] = 8'h15;
mem[16'h6E8F] = 8'h85;
mem[16'h6E90] = 8'h24;
mem[16'h6E91] = 8'hA5;
mem[16'h6E92] = 8'h74;
mem[16'h6E93] = 8'h20;
mem[16'h6E94] = 8'hDA;
mem[16'h6E95] = 8'hFD;
mem[16'h6E96] = 8'h60;
mem[16'h6E97] = 8'hA9;
mem[16'h6E98] = 8'h0C;
mem[16'h6E99] = 8'h85;
mem[16'h6E9A] = 8'h25;
mem[16'h6E9B] = 8'hA9;
mem[16'h6E9C] = 8'h0F;
mem[16'h6E9D] = 8'h85;
mem[16'h6E9E] = 8'h24;
mem[16'h6E9F] = 8'hA9;
mem[16'h6EA0] = 8'hF1;
mem[16'h6EA1] = 8'h85;
mem[16'h6EA2] = 8'h59;
mem[16'h6EA3] = 8'hA9;
mem[16'h6EA4] = 8'h6E;
mem[16'h6EA5] = 8'h85;
mem[16'h6EA6] = 8'h5A;
mem[16'h6EA7] = 8'h20;
mem[16'h6EA8] = 8'hD5;
mem[16'h6EA9] = 8'h67;
mem[16'h6EAA] = 8'hA9;
mem[16'h6EAB] = 8'h0C;
mem[16'h6EAC] = 8'h85;
mem[16'h6EAD] = 8'h25;
mem[16'h6EAE] = 8'hA9;
mem[16'h6EAF] = 8'h15;
mem[16'h6EB0] = 8'h85;
mem[16'h6EB1] = 8'h24;
mem[16'h6EB2] = 8'hA5;
mem[16'h6EB3] = 8'h74;
mem[16'h6EB4] = 8'h20;
mem[16'h6EB5] = 8'hDA;
mem[16'h6EB6] = 8'hFD;
mem[16'h6EB7] = 8'hA9;
mem[16'h6EB8] = 8'h5B;
mem[16'h6EB9] = 8'h8D;
mem[16'h6EBA] = 8'hA1;
mem[16'h6EBB] = 8'h55;
mem[16'h6EBC] = 8'hA9;
mem[16'h6EBD] = 8'h5E;
mem[16'h6EBE] = 8'h8D;
mem[16'h6EBF] = 8'hA2;
mem[16'h6EC0] = 8'h55;
mem[16'h6EC1] = 8'h20;
mem[16'h6EC2] = 8'h51;
mem[16'h6EC3] = 8'h55;
mem[16'h6EC4] = 8'hA9;
mem[16'h6EC5] = 8'h63;
mem[16'h6EC6] = 8'h8D;
mem[16'h6EC7] = 8'hA2;
mem[16'h6EC8] = 8'h55;
mem[16'h6EC9] = 8'h20;
mem[16'h6ECA] = 8'h51;
mem[16'h6ECB] = 8'h55;
mem[16'h6ECC] = 8'hAD;
mem[16'h6ECD] = 8'hA1;
mem[16'h6ECE] = 8'h55;
mem[16'h6ECF] = 8'h18;
mem[16'h6ED0] = 8'h69;
mem[16'h6ED1] = 8'h08;
mem[16'h6ED2] = 8'h8D;
mem[16'h6ED3] = 8'hA1;
mem[16'h6ED4] = 8'h55;
mem[16'h6ED5] = 8'h8D;
mem[16'h6ED6] = 8'hA1;
mem[16'h6ED7] = 8'h55;
mem[16'h6ED8] = 8'hC9;
mem[16'h6ED9] = 8'hB0;
mem[16'h6EDA] = 8'h90;
mem[16'h6EDB] = 8'hE0;
mem[16'h6EDC] = 8'hA9;
mem[16'h6EDD] = 8'h00;
mem[16'h6EDE] = 8'h85;
mem[16'h6EDF] = 8'h70;
mem[16'h6EE0] = 8'hAD;
mem[16'h6EE1] = 8'hC0;
mem[16'h6EE2] = 8'h62;
mem[16'h6EE3] = 8'hF0;
mem[16'h6EE4] = 8'h03;
mem[16'h6EE5] = 8'h20;
mem[16'h6EE6] = 8'hF8;
mem[16'h6EE7] = 8'h62;
mem[16'h6EE8] = 8'hAD;
mem[16'h6EE9] = 8'hC2;
mem[16'h6EEA] = 8'h62;
mem[16'h6EEB] = 8'hF0;
mem[16'h6EEC] = 8'h03;
mem[16'h6EED] = 8'h20;
mem[16'h6EEE] = 8'hC4;
mem[16'h6EEF] = 8'h62;
mem[16'h6EF0] = 8'h60;
mem[16'h6EF1] = 8'hA0;
mem[16'h6EF2] = 8'hD4;
mem[16'h6EF3] = 8'hC9;
mem[16'h6EF4] = 8'hCD;
mem[16'h6EF5] = 8'hC5;
mem[16'h6EF6] = 8'hA0;
mem[16'h6EF7] = 8'h00;
mem[16'h6EF8] = 8'hAD;
mem[16'h6EF9] = 8'h91;
mem[16'h6EFA] = 8'h6F;
mem[16'h6EFB] = 8'h85;
mem[16'h6EFC] = 8'h57;
mem[16'h6EFD] = 8'hA9;
mem[16'h6EFE] = 8'h0A;
mem[16'h6EFF] = 8'h85;
mem[16'h6F00] = 8'h56;
mem[16'h6F01] = 8'hA9;
mem[16'h6F02] = 8'h0A;
mem[16'h6F03] = 8'h8D;
mem[16'h6F04] = 8'hA5;
mem[16'h6F05] = 8'h71;
mem[16'h6F06] = 8'h20;
mem[16'h6F07] = 8'h5E;
mem[16'h6F08] = 8'h71;
mem[16'h6F09] = 8'hA9;
mem[16'h6F0A] = 8'h0A;
mem[16'h6F0B] = 8'h85;
mem[16'h6F0C] = 8'h56;
mem[16'h6F0D] = 8'hA5;
mem[16'h6F0E] = 8'h57;
mem[16'h6F0F] = 8'h18;
mem[16'h6F10] = 8'h69;
mem[16'h6F11] = 8'h08;
mem[16'h6F12] = 8'h85;
mem[16'h6F13] = 8'h57;
mem[16'h6F14] = 8'h20;
mem[16'h6F15] = 8'h5E;
mem[16'h6F16] = 8'h71;
mem[16'h6F17] = 8'hA9;
mem[16'h6F18] = 8'h0A;
mem[16'h6F19] = 8'h85;
mem[16'h6F1A] = 8'h56;
mem[16'h6F1B] = 8'hA5;
mem[16'h6F1C] = 8'h57;
mem[16'h6F1D] = 8'h18;
mem[16'h6F1E] = 8'h69;
mem[16'h6F1F] = 8'h08;
mem[16'h6F20] = 8'h85;
mem[16'h6F21] = 8'h57;
mem[16'h6F22] = 8'h20;
mem[16'h6F23] = 8'h5E;
mem[16'h6F24] = 8'h71;
mem[16'h6F25] = 8'hA9;
mem[16'h6F26] = 8'h0A;
mem[16'h6F27] = 8'h85;
mem[16'h6F28] = 8'h56;
mem[16'h6F29] = 8'hAD;
mem[16'h6F2A] = 8'h91;
mem[16'h6F2B] = 8'h6F;
mem[16'h6F2C] = 8'h85;
mem[16'h6F2D] = 8'h57;
mem[16'h6F2E] = 8'hA9;
mem[16'h6F2F] = 8'h1B;
mem[16'h6F30] = 8'h8D;
mem[16'h6F31] = 8'h7F;
mem[16'h6F32] = 8'h68;
mem[16'h6F33] = 8'h20;
mem[16'h6F34] = 8'hE6;
mem[16'h6F35] = 8'h67;
mem[16'h6F36] = 8'h60;
mem[16'h6F37] = 8'hA9;
mem[16'h6F38] = 8'h0A;
mem[16'h6F39] = 8'h85;
mem[16'h6F3A] = 8'h56;
mem[16'h6F3B] = 8'hAD;
mem[16'h6F3C] = 8'h91;
mem[16'h6F3D] = 8'h6F;
mem[16'h6F3E] = 8'h85;
mem[16'h6F3F] = 8'h57;
mem[16'h6F40] = 8'hA9;
mem[16'h6F41] = 8'h1B;
mem[16'h6F42] = 8'h8D;
mem[16'h6F43] = 8'h7F;
mem[16'h6F44] = 8'h68;
mem[16'h6F45] = 8'h20;
mem[16'h6F46] = 8'hE6;
mem[16'h6F47] = 8'h67;
mem[16'h6F48] = 8'hA9;
mem[16'h6F49] = 8'h0A;
mem[16'h6F4A] = 8'h8D;
mem[16'h6F4B] = 8'hA2;
mem[16'h6F4C] = 8'h55;
mem[16'h6F4D] = 8'hAD;
mem[16'h6F4E] = 8'h91;
mem[16'h6F4F] = 8'h6F;
mem[16'h6F50] = 8'h8D;
mem[16'h6F51] = 8'hA1;
mem[16'h6F52] = 8'h55;
mem[16'h6F53] = 8'h20;
mem[16'h6F54] = 8'h51;
mem[16'h6F55] = 8'h55;
mem[16'h6F56] = 8'hA9;
mem[16'h6F57] = 8'h0F;
mem[16'h6F58] = 8'h8D;
mem[16'h6F59] = 8'hA2;
mem[16'h6F5A] = 8'h55;
mem[16'h6F5B] = 8'h20;
mem[16'h6F5C] = 8'h51;
mem[16'h6F5D] = 8'h55;
mem[16'h6F5E] = 8'hA9;
mem[16'h6F5F] = 8'h0A;
mem[16'h6F60] = 8'h8D;
mem[16'h6F61] = 8'hA2;
mem[16'h6F62] = 8'h55;
mem[16'h6F63] = 8'hAD;
mem[16'h6F64] = 8'hA1;
mem[16'h6F65] = 8'h55;
mem[16'h6F66] = 8'h18;
mem[16'h6F67] = 8'h69;
mem[16'h6F68] = 8'h08;
mem[16'h6F69] = 8'h8D;
mem[16'h6F6A] = 8'hA1;
mem[16'h6F6B] = 8'h55;
mem[16'h6F6C] = 8'h20;
mem[16'h6F6D] = 8'h51;
mem[16'h6F6E] = 8'h55;
mem[16'h6F6F] = 8'hA9;
mem[16'h6F70] = 8'h0F;
mem[16'h6F71] = 8'h8D;
mem[16'h6F72] = 8'hA2;
mem[16'h6F73] = 8'h55;
mem[16'h6F74] = 8'h20;
mem[16'h6F75] = 8'h51;
mem[16'h6F76] = 8'h55;
mem[16'h6F77] = 8'hA9;
mem[16'h6F78] = 8'h0A;
mem[16'h6F79] = 8'h8D;
mem[16'h6F7A] = 8'hA2;
mem[16'h6F7B] = 8'h55;
mem[16'h6F7C] = 8'hAD;
mem[16'h6F7D] = 8'hA1;
mem[16'h6F7E] = 8'h55;
mem[16'h6F7F] = 8'h18;
mem[16'h6F80] = 8'h69;
mem[16'h6F81] = 8'h08;
mem[16'h6F82] = 8'h8D;
mem[16'h6F83] = 8'hA1;
mem[16'h6F84] = 8'h55;
mem[16'h6F85] = 8'h20;
mem[16'h6F86] = 8'h51;
mem[16'h6F87] = 8'h55;
mem[16'h6F88] = 8'hA9;
mem[16'h6F89] = 8'h0F;
mem[16'h6F8A] = 8'h8D;
mem[16'h6F8B] = 8'hA2;
mem[16'h6F8C] = 8'h55;
mem[16'h6F8D] = 8'h20;
mem[16'h6F8E] = 8'h51;
mem[16'h6F8F] = 8'h55;
mem[16'h6F90] = 8'h60;
mem[16'h6F91] = 8'h00;
mem[16'h6F92] = 8'h00;
mem[16'h6F93] = 8'h00;
mem[16'h6F94] = 8'h00;
mem[16'h6F95] = 8'h30;
mem[16'h6F96] = 8'h18;
mem[16'h6F97] = 8'h0C;
mem[16'h6F98] = 8'h48;
mem[16'h6F99] = 8'h24;
mem[16'h6F9A] = 8'h12;
mem[16'h6F9B] = 8'h40;
mem[16'h6F9C] = 8'h24;
mem[16'h6F9D] = 8'h12;
mem[16'h6F9E] = 8'h20;
mem[16'h6F9F] = 8'h24;
mem[16'h6FA0] = 8'h12;
mem[16'h6FA1] = 8'h18;
mem[16'h6FA2] = 8'h24;
mem[16'h6FA3] = 8'h12;
mem[16'h6FA4] = 8'h08;
mem[16'h6FA5] = 8'h24;
mem[16'h6FA6] = 8'h12;
mem[16'h6FA7] = 8'h78;
mem[16'h6FA8] = 8'h18;
mem[16'h6FA9] = 8'h0C;
mem[16'h6FAA] = 8'h00;
mem[16'h6FAB] = 8'h00;
mem[16'h6FAC] = 8'h00;
mem[16'h6FAD] = 8'h00;
mem[16'h6FAE] = 8'h00;
mem[16'h6FAF] = 8'h00;
mem[16'h6FB0] = 8'h24;
mem[16'h6FB1] = 8'h18;
mem[16'h6FB2] = 8'h0C;
mem[16'h6FB3] = 8'h24;
mem[16'h6FB4] = 8'h24;
mem[16'h6FB5] = 8'h12;
mem[16'h6FB6] = 8'h24;
mem[16'h6FB7] = 8'h24;
mem[16'h6FB8] = 8'h12;
mem[16'h6FB9] = 8'h7C;
mem[16'h6FBA] = 8'h24;
mem[16'h6FBB] = 8'h12;
mem[16'h6FBC] = 8'h20;
mem[16'h6FBD] = 8'h24;
mem[16'h6FBE] = 8'h12;
mem[16'h6FBF] = 8'h20;
mem[16'h6FC0] = 8'h24;
mem[16'h6FC1] = 8'h12;
mem[16'h6FC2] = 8'h20;
mem[16'h6FC3] = 8'h18;
mem[16'h6FC4] = 8'h0C;
mem[16'h6FC5] = 8'h00;
mem[16'h6FC6] = 8'h00;
mem[16'h6FC7] = 8'h00;
mem[16'h6FC8] = 8'hA9;
mem[16'h6FC9] = 8'h41;
mem[16'h6FCA] = 8'h85;
mem[16'h6FCB] = 8'h79;
mem[16'h6FCC] = 8'hA9;
mem[16'h6FCD] = 8'h83;
mem[16'h6FCE] = 8'h85;
mem[16'h6FCF] = 8'h7A;
mem[16'h6FD0] = 8'hA9;
mem[16'h6FD1] = 8'h7E;
mem[16'h6FD2] = 8'h85;
mem[16'h6FD3] = 8'h7B;
mem[16'h6FD4] = 8'hA9;
mem[16'h6FD5] = 8'h83;
mem[16'h6FD6] = 8'h85;
mem[16'h6FD7] = 8'h7C;
mem[16'h6FD8] = 8'h20;
mem[16'h6FD9] = 8'hA2;
mem[16'h6FDA] = 8'h82;
mem[16'h6FDB] = 8'h60;
mem[16'h6FDC] = 8'hAD;
mem[16'h6FDD] = 8'h00;
mem[16'h6FDE] = 8'hC0;
mem[16'h6FDF] = 8'hC9;
mem[16'h6FE0] = 8'h9B;
mem[16'h6FE1] = 8'hD0;
mem[16'h6FE2] = 8'h0D;
mem[16'h6FE3] = 8'hAD;
mem[16'h6FE4] = 8'h10;
mem[16'h6FE5] = 8'hC0;
mem[16'h6FE6] = 8'hAD;
mem[16'h6FE7] = 8'h00;
mem[16'h6FE8] = 8'hC0;
mem[16'h6FE9] = 8'hC9;
mem[16'h6FEA] = 8'h9B;
mem[16'h6FEB] = 8'hD0;
mem[16'h6FEC] = 8'hF9;
mem[16'h6FED] = 8'hAD;
mem[16'h6FEE] = 8'h10;
mem[16'h6FEF] = 8'hC0;
mem[16'h6FF0] = 8'h60;
mem[16'h6FF1] = 8'hCE;
mem[16'h6FF2] = 8'h22;
mem[16'h6FF3] = 8'h70;
mem[16'h6FF4] = 8'hAE;
mem[16'h6FF5] = 8'h22;
mem[16'h6FF6] = 8'h70;
mem[16'h6FF7] = 8'hBD;
mem[16'h6FF8] = 8'h76;
mem[16'h6FF9] = 8'h41;
mem[16'h6FFA] = 8'h1D;
mem[16'h6FFB] = 8'h2A;
mem[16'h6FFC] = 8'h61;
mem[16'h6FFD] = 8'h45;
mem[16'h6FFE] = 8'h73;
mem[16'h6FFF] = 8'h29;
mem[16'h7000] = 8'h03;
mem[16'h7001] = 8'hD0;
mem[16'h7002] = 8'h1E;
mem[16'h7003] = 8'hA5;
mem[16'h7004] = 8'h73;
mem[16'h7005] = 8'hC9;
mem[16'h7006] = 8'h01;
mem[16'h7007] = 8'hD0;
mem[16'h7008] = 8'h03;
mem[16'h7009] = 8'h20;
mem[16'h700A] = 8'hFF;
mem[16'h700B] = 8'h55;
mem[16'h700C] = 8'hA5;
mem[16'h700D] = 8'h73;
mem[16'h700E] = 8'hC9;
mem[16'h700F] = 8'h02;
mem[16'h7010] = 8'hD0;
mem[16'h7011] = 8'h07;
mem[16'h7012] = 8'h20;
mem[16'h7013] = 8'h28;
mem[16'h7014] = 8'h5C;
mem[16'h7015] = 8'h20;
mem[16'h7016] = 8'h87;
mem[16'h7017] = 8'h58;
mem[16'h7018] = 8'h60;
mem[16'h7019] = 8'hA5;
mem[16'h701A] = 8'h73;
mem[16'h701B] = 8'h20;
mem[16'h701C] = 8'h62;
mem[16'h701D] = 8'h5C;
mem[16'h701E] = 8'h20;
mem[16'h701F] = 8'h43;
mem[16'h7020] = 8'h57;
mem[16'h7021] = 8'h60;
mem[16'h7022] = 8'h20;
mem[16'h7023] = 8'h20;
mem[16'h7024] = 8'h42;
mem[16'h7025] = 8'h65;
mem[16'h7026] = 8'h20;
mem[16'h7027] = 8'h2F;
mem[16'h7028] = 8'h65;
mem[16'h7029] = 8'hAD;
mem[16'h702A] = 8'h10;
mem[16'h702B] = 8'hC0;
mem[16'h702C] = 8'hA9;
mem[16'h702D] = 8'hD4;
mem[16'h702E] = 8'h85;
mem[16'h702F] = 8'h59;
mem[16'h7030] = 8'hA9;
mem[16'h7031] = 8'h70;
mem[16'h7032] = 8'h85;
mem[16'h7033] = 8'h5A;
mem[16'h7034] = 8'hA9;
mem[16'h7035] = 8'h0A;
mem[16'h7036] = 8'h85;
mem[16'h7037] = 8'h24;
mem[16'h7038] = 8'hA9;
mem[16'h7039] = 8'h01;
mem[16'h703A] = 8'h85;
mem[16'h703B] = 8'h25;
mem[16'h703C] = 8'h20;
mem[16'h703D] = 8'hD5;
mem[16'h703E] = 8'h67;
mem[16'h703F] = 8'hA9;
mem[16'h7040] = 8'hE2;
mem[16'h7041] = 8'h85;
mem[16'h7042] = 8'h59;
mem[16'h7043] = 8'hA9;
mem[16'h7044] = 8'h70;
mem[16'h7045] = 8'h85;
mem[16'h7046] = 8'h5A;
mem[16'h7047] = 8'hA9;
mem[16'h7048] = 8'h08;
mem[16'h7049] = 8'h85;
mem[16'h704A] = 8'h24;
mem[16'h704B] = 8'hA9;
mem[16'h704C] = 8'h06;
mem[16'h704D] = 8'h85;
mem[16'h704E] = 8'h25;
mem[16'h704F] = 8'h20;
mem[16'h7050] = 8'hD5;
mem[16'h7051] = 8'h67;
mem[16'h7052] = 8'hAD;
mem[16'h7053] = 8'h00;
mem[16'h7054] = 8'hC0;
mem[16'h7055] = 8'h29;
mem[16'h7056] = 8'h80;
mem[16'h7057] = 8'hF0;
mem[16'h7058] = 8'hF9;
mem[16'h7059] = 8'hAD;
mem[16'h705A] = 8'h00;
mem[16'h705B] = 8'hC0;
mem[16'h705C] = 8'h85;
mem[16'h705D] = 8'h7D;
mem[16'h705E] = 8'h20;
mem[16'h705F] = 8'hED;
mem[16'h7060] = 8'hFD;
mem[16'h7061] = 8'hAD;
mem[16'h7062] = 8'h10;
mem[16'h7063] = 8'hC0;
mem[16'h7064] = 8'hA9;
mem[16'h7065] = 8'hFA;
mem[16'h7066] = 8'h85;
mem[16'h7067] = 8'h59;
mem[16'h7068] = 8'hA9;
mem[16'h7069] = 8'h70;
mem[16'h706A] = 8'h85;
mem[16'h706B] = 8'h5A;
mem[16'h706C] = 8'hA9;
mem[16'h706D] = 8'h08;
mem[16'h706E] = 8'h85;
mem[16'h706F] = 8'h24;
mem[16'h7070] = 8'hA9;
mem[16'h7071] = 8'h08;
mem[16'h7072] = 8'h85;
mem[16'h7073] = 8'h25;
mem[16'h7074] = 8'h20;
mem[16'h7075] = 8'hD5;
mem[16'h7076] = 8'h67;
mem[16'h7077] = 8'hAD;
mem[16'h7078] = 8'h00;
mem[16'h7079] = 8'hC0;
mem[16'h707A] = 8'h29;
mem[16'h707B] = 8'h80;
mem[16'h707C] = 8'hF0;
mem[16'h707D] = 8'hF9;
mem[16'h707E] = 8'hAD;
mem[16'h707F] = 8'h00;
mem[16'h7080] = 8'hC0;
mem[16'h7081] = 8'h85;
mem[16'h7082] = 8'h7E;
mem[16'h7083] = 8'h20;
mem[16'h7084] = 8'hED;
mem[16'h7085] = 8'hFD;
mem[16'h7086] = 8'hAD;
mem[16'h7087] = 8'h10;
mem[16'h7088] = 8'hC0;
mem[16'h7089] = 8'hA9;
mem[16'h708A] = 8'h14;
mem[16'h708B] = 8'h85;
mem[16'h708C] = 8'h59;
mem[16'h708D] = 8'hA9;
mem[16'h708E] = 8'h71;
mem[16'h708F] = 8'h85;
mem[16'h7090] = 8'h5A;
mem[16'h7091] = 8'hA9;
mem[16'h7092] = 8'h08;
mem[16'h7093] = 8'h85;
mem[16'h7094] = 8'h24;
mem[16'h7095] = 8'hA9;
mem[16'h7096] = 8'h0A;
mem[16'h7097] = 8'h85;
mem[16'h7098] = 8'h25;
mem[16'h7099] = 8'h20;
mem[16'h709A] = 8'hD5;
mem[16'h709B] = 8'h67;
mem[16'h709C] = 8'hAD;
mem[16'h709D] = 8'h00;
mem[16'h709E] = 8'hC0;
mem[16'h709F] = 8'h29;
mem[16'h70A0] = 8'h80;
mem[16'h70A1] = 8'hF0;
mem[16'h70A2] = 8'hF9;
mem[16'h70A3] = 8'hAD;
mem[16'h70A4] = 8'h00;
mem[16'h70A5] = 8'hC0;
mem[16'h70A6] = 8'h85;
mem[16'h70A7] = 8'h80;
mem[16'h70A8] = 8'h20;
mem[16'h70A9] = 8'hED;
mem[16'h70AA] = 8'hFD;
mem[16'h70AB] = 8'hAD;
mem[16'h70AC] = 8'h10;
mem[16'h70AD] = 8'hC0;
mem[16'h70AE] = 8'hA9;
mem[16'h70AF] = 8'h2F;
mem[16'h70B0] = 8'h85;
mem[16'h70B1] = 8'h59;
mem[16'h70B2] = 8'hA9;
mem[16'h70B3] = 8'h71;
mem[16'h70B4] = 8'h85;
mem[16'h70B5] = 8'h5A;
mem[16'h70B6] = 8'hA9;
mem[16'h70B7] = 8'h08;
mem[16'h70B8] = 8'h85;
mem[16'h70B9] = 8'h24;
mem[16'h70BA] = 8'hA9;
mem[16'h70BB] = 8'h0C;
mem[16'h70BC] = 8'h85;
mem[16'h70BD] = 8'h25;
mem[16'h70BE] = 8'h20;
mem[16'h70BF] = 8'hD5;
mem[16'h70C0] = 8'h67;
mem[16'h70C1] = 8'hAD;
mem[16'h70C2] = 8'h00;
mem[16'h70C3] = 8'hC0;
mem[16'h70C4] = 8'h29;
mem[16'h70C5] = 8'h80;
mem[16'h70C6] = 8'hF0;
mem[16'h70C7] = 8'hF9;
mem[16'h70C8] = 8'hAD;
mem[16'h70C9] = 8'h00;
mem[16'h70CA] = 8'hC0;
mem[16'h70CB] = 8'h85;
mem[16'h70CC] = 8'h7F;
mem[16'h70CD] = 8'h20;
mem[16'h70CE] = 8'hED;
mem[16'h70CF] = 8'hFD;
mem[16'h70D0] = 8'hAD;
mem[16'h70D1] = 8'h10;
mem[16'h70D2] = 8'hC0;
mem[16'h70D3] = 8'h60;
mem[16'h70D4] = 8'hD2;
mem[16'h70D5] = 8'hC5;
mem[16'h70D6] = 8'hC4;
mem[16'h70D7] = 8'hC5;
mem[16'h70D8] = 8'hC6;
mem[16'h70D9] = 8'hC9;
mem[16'h70DA] = 8'hCE;
mem[16'h70DB] = 8'hC5;
mem[16'h70DC] = 8'hA0;
mem[16'h70DD] = 8'hCB;
mem[16'h70DE] = 8'hC5;
mem[16'h70DF] = 8'hD9;
mem[16'h70E0] = 8'hD3;
mem[16'h70E1] = 8'h00;
mem[16'h70E2] = 8'hD4;
mem[16'h70E3] = 8'hD9;
mem[16'h70E4] = 8'hD0;
mem[16'h70E5] = 8'hC5;
mem[16'h70E6] = 8'hA0;
mem[16'h70E7] = 8'hC9;
mem[16'h70E8] = 8'hCE;
mem[16'h70E9] = 8'hA0;
mem[16'h70EA] = 8'hD4;
mem[16'h70EB] = 8'hC8;
mem[16'h70EC] = 8'hC5;
mem[16'h70ED] = 8'hA0;
mem[16'h70EE] = 8'hA7;
mem[16'h70EF] = 8'hD5;
mem[16'h70F0] = 8'hD0;
mem[16'h70F1] = 8'hA7;
mem[16'h70F2] = 8'hA0;
mem[16'h70F3] = 8'hCB;
mem[16'h70F4] = 8'hC5;
mem[16'h70F5] = 8'hD9;
mem[16'h70F6] = 8'hA0;
mem[16'h70F7] = 8'hAD;
mem[16'h70F8] = 8'hA0;
mem[16'h70F9] = 8'h00;
mem[16'h70FA] = 8'hD4;
mem[16'h70FB] = 8'hD9;
mem[16'h70FC] = 8'hD0;
mem[16'h70FD] = 8'hC5;
mem[16'h70FE] = 8'hA0;
mem[16'h70FF] = 8'hC9;
mem[16'h7100] = 8'hCE;
mem[16'h7101] = 8'hA0;
mem[16'h7102] = 8'hD4;
mem[16'h7103] = 8'hC8;
mem[16'h7104] = 8'hC5;
mem[16'h7105] = 8'hA0;
mem[16'h7106] = 8'hA7;
mem[16'h7107] = 8'hC4;
mem[16'h7108] = 8'hCF;
mem[16'h7109] = 8'hD7;
mem[16'h710A] = 8'hCE;
mem[16'h710B] = 8'hA7;
mem[16'h710C] = 8'hA0;
mem[16'h710D] = 8'hCB;
mem[16'h710E] = 8'hC5;
mem[16'h710F] = 8'hD9;
mem[16'h7110] = 8'hA0;
mem[16'h7111] = 8'hAD;
mem[16'h7112] = 8'hA0;
mem[16'h7113] = 8'h00;
mem[16'h7114] = 8'hD4;
mem[16'h7115] = 8'hD9;
mem[16'h7116] = 8'hD0;
mem[16'h7117] = 8'hC5;
mem[16'h7118] = 8'hA0;
mem[16'h7119] = 8'hC9;
mem[16'h711A] = 8'hCE;
mem[16'h711B] = 8'hA0;
mem[16'h711C] = 8'hD4;
mem[16'h711D] = 8'hC8;
mem[16'h711E] = 8'hC5;
mem[16'h711F] = 8'hA0;
mem[16'h7120] = 8'hA7;
mem[16'h7121] = 8'hD2;
mem[16'h7122] = 8'hC9;
mem[16'h7123] = 8'hC7;
mem[16'h7124] = 8'hC8;
mem[16'h7125] = 8'hD4;
mem[16'h7126] = 8'hA7;
mem[16'h7127] = 8'hA0;
mem[16'h7128] = 8'hCB;
mem[16'h7129] = 8'hC5;
mem[16'h712A] = 8'hD9;
mem[16'h712B] = 8'hA0;
mem[16'h712C] = 8'hAD;
mem[16'h712D] = 8'hA0;
mem[16'h712E] = 8'h00;
mem[16'h712F] = 8'hD4;
mem[16'h7130] = 8'hD9;
mem[16'h7131] = 8'hD0;
mem[16'h7132] = 8'hC5;
mem[16'h7133] = 8'hA0;
mem[16'h7134] = 8'hC9;
mem[16'h7135] = 8'hCE;
mem[16'h7136] = 8'hA0;
mem[16'h7137] = 8'hD4;
mem[16'h7138] = 8'hC8;
mem[16'h7139] = 8'hC5;
mem[16'h713A] = 8'hA0;
mem[16'h713B] = 8'hA7;
mem[16'h713C] = 8'hCC;
mem[16'h713D] = 8'hC5;
mem[16'h713E] = 8'hC6;
mem[16'h713F] = 8'hD4;
mem[16'h7140] = 8'hA7;
mem[16'h7141] = 8'hA0;
mem[16'h7142] = 8'hCB;
mem[16'h7143] = 8'hC5;
mem[16'h7144] = 8'hD9;
mem[16'h7145] = 8'hA0;
mem[16'h7146] = 8'hAD;
mem[16'h7147] = 8'hA0;
mem[16'h7148] = 8'h00;
mem[16'h7149] = 8'hA9;
mem[16'h714A] = 8'hC1;
mem[16'h714B] = 8'h85;
mem[16'h714C] = 8'h7D;
mem[16'h714D] = 8'hA9;
mem[16'h714E] = 8'hDA;
mem[16'h714F] = 8'h85;
mem[16'h7150] = 8'h7E;
mem[16'h7151] = 8'hA9;
mem[16'h7152] = 8'h88;
mem[16'h7153] = 8'h85;
mem[16'h7154] = 8'h7F;
mem[16'h7155] = 8'hA9;
mem[16'h7156] = 8'h95;
mem[16'h7157] = 8'h85;
mem[16'h7158] = 8'h80;
mem[16'h7159] = 8'hA9;
mem[16'h715A] = 8'h00;
mem[16'h715B] = 8'h85;
mem[16'h715C] = 8'h85;
mem[16'h715D] = 8'h60;
mem[16'h715E] = 8'hA2;
mem[16'h715F] = 8'h00;
mem[16'h7160] = 8'hA4;
mem[16'h7161] = 8'h56;
mem[16'h7162] = 8'hB9;
mem[16'h7163] = 8'hD5;
mem[16'h7164] = 8'h8E;
mem[16'h7165] = 8'h85;
mem[16'h7166] = 8'h59;
mem[16'h7167] = 8'hB9;
mem[16'h7168] = 8'h95;
mem[16'h7169] = 8'h8F;
mem[16'h716A] = 8'h85;
mem[16'h716B] = 8'h5A;
mem[16'h716C] = 8'hA4;
mem[16'h716D] = 8'h57;
mem[16'h716E] = 8'hB9;
mem[16'h716F] = 8'h3E;
mem[16'h7170] = 8'h8C;
mem[16'h7171] = 8'h85;
mem[16'h7172] = 8'h5C;
mem[16'h7173] = 8'hB9;
mem[16'h7174] = 8'h56;
mem[16'h7175] = 8'h8D;
mem[16'h7176] = 8'hA8;
mem[16'h7177] = 8'hA9;
mem[16'h7178] = 8'h00;
mem[16'h7179] = 8'h85;
mem[16'h717A] = 8'h6D;
mem[16'h717B] = 8'h85;
mem[16'h717C] = 8'h66;
mem[16'h717D] = 8'hA9;
mem[16'h717E] = 8'hFF;
mem[16'h717F] = 8'h85;
mem[16'h7180] = 8'h6A;
mem[16'h7181] = 8'hA5;
mem[16'h7182] = 8'h5C;
mem[16'h7183] = 8'hC9;
mem[16'h7184] = 8'h01;
mem[16'h7185] = 8'hF0;
mem[16'h7186] = 8'h14;
mem[16'h7187] = 8'h38;
mem[16'h7188] = 8'h66;
mem[16'h7189] = 8'h66;
mem[16'h718A] = 8'h66;
mem[16'h718B] = 8'h6A;
mem[16'h718C] = 8'h06;
mem[16'h718D] = 8'h5C;
mem[16'h718E] = 8'h24;
mem[16'h718F] = 8'h5C;
mem[16'h7190] = 8'h10;
mem[16'h7191] = 8'hF5;
mem[16'h7192] = 8'h46;
mem[16'h7193] = 8'h6A;
mem[16'h7194] = 8'hA5;
mem[16'h7195] = 8'h6A;
mem[16'h7196] = 8'h31;
mem[16'h7197] = 8'h59;
mem[16'h7198] = 8'h91;
mem[16'h7199] = 8'h59;
mem[16'h719A] = 8'hC8;
mem[16'h719B] = 8'hA5;
mem[16'h719C] = 8'h66;
mem[16'h719D] = 8'h31;
mem[16'h719E] = 8'h59;
mem[16'h719F] = 8'h91;
mem[16'h71A0] = 8'h59;
mem[16'h71A1] = 8'hE6;
mem[16'h71A2] = 8'h56;
mem[16'h71A3] = 8'hE8;
mem[16'h71A4] = 8'hE0;
mem[16'h71A5] = 8'h07;
mem[16'h71A6] = 8'hB0;
mem[16'h71A7] = 8'h03;
mem[16'h71A8] = 8'h4C;
mem[16'h71A9] = 8'h60;
mem[16'h71AA] = 8'h71;
mem[16'h71AB] = 8'h60;
mem[16'h71AC] = 8'hA2;
mem[16'h71AD] = 8'h00;
mem[16'h71AE] = 8'hA4;
mem[16'h71AF] = 8'h56;
mem[16'h71B0] = 8'hC0;
mem[16'h71B1] = 8'hC0;
mem[16'h71B2] = 8'h90;
mem[16'h71B3] = 8'h06;
mem[16'h71B4] = 8'h20;
mem[16'h71B5] = 8'hDD;
mem[16'h71B6] = 8'hFB;
mem[16'h71B7] = 8'h4C;
mem[16'h71B8] = 8'hF3;
mem[16'h71B9] = 8'h71;
mem[16'h71BA] = 8'hB9;
mem[16'h71BB] = 8'hD5;
mem[16'h71BC] = 8'h8E;
mem[16'h71BD] = 8'h85;
mem[16'h71BE] = 8'h59;
mem[16'h71BF] = 8'hB9;
mem[16'h71C0] = 8'h95;
mem[16'h71C1] = 8'h8F;
mem[16'h71C2] = 8'h85;
mem[16'h71C3] = 8'h5A;
mem[16'h71C4] = 8'hA4;
mem[16'h71C5] = 8'h57;
mem[16'h71C6] = 8'hB9;
mem[16'h71C7] = 8'h56;
mem[16'h71C8] = 8'h8D;
mem[16'h71C9] = 8'hA8;
mem[16'h71CA] = 8'hBD;
mem[16'h71CB] = 8'h8D;
mem[16'h71CC] = 8'h80;
mem[16'h71CD] = 8'h29;
mem[16'h71CE] = 8'h80;
mem[16'h71CF] = 8'h85;
mem[16'h71D0] = 8'h6D;
mem[16'h71D1] = 8'hBD;
mem[16'h71D2] = 8'h8D;
mem[16'h71D3] = 8'h80;
mem[16'h71D4] = 8'h29;
mem[16'h71D5] = 8'h7F;
mem[16'h71D6] = 8'h51;
mem[16'h71D7] = 8'h59;
mem[16'h71D8] = 8'h05;
mem[16'h71D9] = 8'h6D;
mem[16'h71DA] = 8'h91;
mem[16'h71DB] = 8'h59;
mem[16'h71DC] = 8'hE8;
mem[16'h71DD] = 8'hC8;
mem[16'h71DE] = 8'hBD;
mem[16'h71DF] = 8'h8D;
mem[16'h71E0] = 8'h80;
mem[16'h71E1] = 8'h29;
mem[16'h71E2] = 8'h7F;
mem[16'h71E3] = 8'h51;
mem[16'h71E4] = 8'h59;
mem[16'h71E5] = 8'h05;
mem[16'h71E6] = 8'h6D;
mem[16'h71E7] = 8'h91;
mem[16'h71E8] = 8'h59;
mem[16'h71E9] = 8'hE6;
mem[16'h71EA] = 8'h56;
mem[16'h71EB] = 8'hE8;
mem[16'h71EC] = 8'hE0;
mem[16'h71ED] = 8'h12;
mem[16'h71EE] = 8'hB0;
mem[16'h71EF] = 8'h03;
mem[16'h71F0] = 8'h4C;
mem[16'h71F1] = 8'hAE;
mem[16'h71F2] = 8'h71;
mem[16'h71F3] = 8'h60;
mem[16'h71F4] = 8'h8D;
mem[16'h71F5] = 8'hCB;
mem[16'h71F6] = 8'h71;
mem[16'h71F7] = 8'h8D;
mem[16'h71F8] = 8'hD2;
mem[16'h71F9] = 8'h71;
mem[16'h71FA] = 8'h8D;
mem[16'h71FB] = 8'hDF;
mem[16'h71FC] = 8'h71;
mem[16'h71FD] = 8'h8C;
mem[16'h71FE] = 8'hCC;
mem[16'h71FF] = 8'h71;
mem[16'h7200] = 8'h8C;
mem[16'h7201] = 8'hD3;
mem[16'h7202] = 8'h71;
mem[16'h7203] = 8'h8C;
mem[16'h7204] = 8'hE0;
mem[16'h7205] = 8'h71;
mem[16'h7206] = 8'h60;
mem[16'h7207] = 8'hC0;
mem[16'h7208] = 8'h5B;
mem[16'h7209] = 8'h03;
mem[16'h720A] = 8'hC0;
mem[16'h720B] = 8'h5B;
mem[16'h720C] = 8'h53;
mem[16'h720D] = 8'hC0;
mem[16'h720E] = 8'h00;
mem[16'h720F] = 8'h2C;
mem[16'h7210] = 8'hC0;
mem[16'h7211] = 8'h00;
mem[16'h7212] = 8'h32;
mem[16'h7213] = 8'hC0;
mem[16'h7214] = 8'h00;
mem[16'h7215] = 8'h2C;
mem[16'h7216] = 8'hC0;
mem[16'h7217] = 8'h00;
mem[16'h7218] = 8'h32;
mem[16'h7219] = 8'hC0;
mem[16'h721A] = 8'h00;
mem[16'h721B] = 8'h2C;
mem[16'h721C] = 8'hC0;
mem[16'h721D] = 8'h5B;
mem[16'h721E] = 8'h53;
mem[16'h721F] = 8'hC0;
mem[16'h7220] = 8'h5B;
mem[16'h7221] = 8'h03;
mem[16'h7222] = 8'hE0;
mem[16'h7223] = 8'h6D;
mem[16'h7224] = 8'h01;
mem[16'h7225] = 8'hE0;
mem[16'h7226] = 8'h6D;
mem[16'h7227] = 8'h29;
mem[16'h7228] = 8'hA0;
mem[16'h7229] = 8'h00;
mem[16'h722A] = 8'h16;
mem[16'h722B] = 8'hA0;
mem[16'h722C] = 8'h00;
mem[16'h722D] = 8'h19;
mem[16'h722E] = 8'hA0;
mem[16'h722F] = 8'h00;
mem[16'h7230] = 8'h16;
mem[16'h7231] = 8'hA0;
mem[16'h7232] = 8'h00;
mem[16'h7233] = 8'h19;
mem[16'h7234] = 8'hA0;
mem[16'h7235] = 8'h00;
mem[16'h7236] = 8'h16;
mem[16'h7237] = 8'hE0;
mem[16'h7238] = 8'h6D;
mem[16'h7239] = 8'h29;
mem[16'h723A] = 8'hE0;
mem[16'h723B] = 8'h6D;
mem[16'h723C] = 8'h01;
mem[16'h723D] = 8'hF0;
mem[16'h723E] = 8'h76;
mem[16'h723F] = 8'h00;
mem[16'h7240] = 8'hF0;
mem[16'h7241] = 8'h76;
mem[16'h7242] = 8'h14;
mem[16'h7243] = 8'h90;
mem[16'h7244] = 8'h00;
mem[16'h7245] = 8'h0B;
mem[16'h7246] = 8'h90;
mem[16'h7247] = 8'h40;
mem[16'h7248] = 8'h0C;
mem[16'h7249] = 8'h90;
mem[16'h724A] = 8'h00;
mem[16'h724B] = 8'h0B;
mem[16'h724C] = 8'h90;
mem[16'h724D] = 8'h40;
mem[16'h724E] = 8'h0C;
mem[16'h724F] = 8'h90;
mem[16'h7250] = 8'h00;
mem[16'h7251] = 8'h0B;
mem[16'h7252] = 8'hF0;
mem[16'h7253] = 8'h76;
mem[16'h7254] = 8'h14;
mem[16'h7255] = 8'hF0;
mem[16'h7256] = 8'h76;
mem[16'h7257] = 8'h00;
mem[16'h7258] = 8'hB8;
mem[16'h7259] = 8'h3B;
mem[16'h725A] = 8'h00;
mem[16'h725B] = 8'hB8;
mem[16'h725C] = 8'h3B;
mem[16'h725D] = 8'h0A;
mem[16'h725E] = 8'h88;
mem[16'h725F] = 8'h40;
mem[16'h7260] = 8'h05;
mem[16'h7261] = 8'h88;
mem[16'h7262] = 8'h20;
mem[16'h7263] = 8'h06;
mem[16'h7264] = 8'h88;
mem[16'h7265] = 8'h40;
mem[16'h7266] = 8'h05;
mem[16'h7267] = 8'h88;
mem[16'h7268] = 8'h20;
mem[16'h7269] = 8'h06;
mem[16'h726A] = 8'h88;
mem[16'h726B] = 8'h40;
mem[16'h726C] = 8'h05;
mem[16'h726D] = 8'hB8;
mem[16'h726E] = 8'h3B;
mem[16'h726F] = 8'h0A;
mem[16'h7270] = 8'hB8;
mem[16'h7271] = 8'h3B;
mem[16'h7272] = 8'h00;
mem[16'h7273] = 8'hDC;
mem[16'h7274] = 8'h1D;
mem[16'h7275] = 8'h00;
mem[16'h7276] = 8'hDC;
mem[16'h7277] = 8'h1D;
mem[16'h7278] = 8'h05;
mem[16'h7279] = 8'h84;
mem[16'h727A] = 8'h60;
mem[16'h727B] = 8'h02;
mem[16'h727C] = 8'h84;
mem[16'h727D] = 8'h10;
mem[16'h727E] = 8'h03;
mem[16'h727F] = 8'h84;
mem[16'h7280] = 8'h60;
mem[16'h7281] = 8'h02;
mem[16'h7282] = 8'h84;
mem[16'h7283] = 8'h10;
mem[16'h7284] = 8'h03;
mem[16'h7285] = 8'h84;
mem[16'h7286] = 8'h60;
mem[16'h7287] = 8'h02;
mem[16'h7288] = 8'hDC;
mem[16'h7289] = 8'h1D;
mem[16'h728A] = 8'h05;
mem[16'h728B] = 8'hDC;
mem[16'h728C] = 8'h1D;
mem[16'h728D] = 8'h00;
mem[16'h728E] = 8'hEE;
mem[16'h728F] = 8'h0E;
mem[16'h7290] = 8'h00;
mem[16'h7291] = 8'hEE;
mem[16'h7292] = 8'h4E;
mem[16'h7293] = 8'h02;
mem[16'h7294] = 8'h82;
mem[16'h7295] = 8'h30;
mem[16'h7296] = 8'h01;
mem[16'h7297] = 8'h82;
mem[16'h7298] = 8'h48;
mem[16'h7299] = 8'h01;
mem[16'h729A] = 8'h82;
mem[16'h729B] = 8'h30;
mem[16'h729C] = 8'h01;
mem[16'h729D] = 8'h82;
mem[16'h729E] = 8'h48;
mem[16'h729F] = 8'h01;
mem[16'h72A0] = 8'h82;
mem[16'h72A1] = 8'h30;
mem[16'h72A2] = 8'h01;
mem[16'h72A3] = 8'hEE;
mem[16'h72A4] = 8'h4E;
mem[16'h72A5] = 8'h02;
mem[16'h72A6] = 8'hEE;
mem[16'h72A7] = 8'h0E;
mem[16'h72A8] = 8'h00;
mem[16'h72A9] = 8'hB7;
mem[16'h72AA] = 8'h07;
mem[16'h72AB] = 8'h00;
mem[16'h72AC] = 8'hB7;
mem[16'h72AD] = 8'h27;
mem[16'h72AE] = 8'h01;
mem[16'h72AF] = 8'h81;
mem[16'h72B0] = 8'h58;
mem[16'h72B1] = 8'h00;
mem[16'h72B2] = 8'h81;
mem[16'h72B3] = 8'h64;
mem[16'h72B4] = 8'h00;
mem[16'h72B5] = 8'h81;
mem[16'h72B6] = 8'h58;
mem[16'h72B7] = 8'h00;
mem[16'h72B8] = 8'h81;
mem[16'h72B9] = 8'h64;
mem[16'h72BA] = 8'h00;
mem[16'h72BB] = 8'h81;
mem[16'h72BC] = 8'h58;
mem[16'h72BD] = 8'h00;
mem[16'h72BE] = 8'hB7;
mem[16'h72BF] = 8'h27;
mem[16'h72C0] = 8'h01;
mem[16'h72C1] = 8'hB7;
mem[16'h72C2] = 8'h07;
mem[16'h72C3] = 8'h00;
mem[16'h72C4] = 8'hA6;
mem[16'h72C5] = 8'h70;
mem[16'h72C6] = 8'hBD;
mem[16'h72C7] = 8'h75;
mem[16'h72C8] = 8'h5B;
mem[16'h72C9] = 8'hD0;
mem[16'h72CA] = 8'h04;
mem[16'h72CB] = 8'h20;
mem[16'h72CC] = 8'hC6;
mem[16'h72CD] = 8'h5E;
mem[16'h72CE] = 8'h60;
mem[16'h72CF] = 8'hC9;
mem[16'h72D0] = 8'h1E;
mem[16'h72D1] = 8'hB0;
mem[16'h72D2] = 8'h04;
mem[16'h72D3] = 8'hC9;
mem[16'h72D4] = 8'h08;
mem[16'h72D5] = 8'hB0;
mem[16'h72D6] = 8'h04;
mem[16'h72D7] = 8'h20;
mem[16'h72D8] = 8'hE8;
mem[16'h72D9] = 8'h72;
mem[16'h72DA] = 8'h60;
mem[16'h72DB] = 8'hC9;
mem[16'h72DC] = 8'h16;
mem[16'h72DD] = 8'hB0;
mem[16'h72DE] = 8'h05;
mem[16'h72DF] = 8'hC9;
mem[16'h72E0] = 8'h0F;
mem[16'h72E1] = 8'h90;
mem[16'h72E2] = 8'h01;
mem[16'h72E3] = 8'h60;
mem[16'h72E4] = 8'h20;
mem[16'h72E5] = 8'hF4;
mem[16'h72E6] = 8'h72;
mem[16'h72E7] = 8'h60;
mem[16'h72E8] = 8'hA9;
mem[16'h72E9] = 8'h16;
mem[16'h72EA] = 8'h8D;
mem[16'h72EB] = 8'h24;
mem[16'h72EC] = 8'h8C;
mem[16'h72ED] = 8'hA9;
mem[16'h72EE] = 8'h6F;
mem[16'h72EF] = 8'hA0;
mem[16'h72F0] = 8'h4F;
mem[16'h72F1] = 8'h4C;
mem[16'h72F2] = 8'hFD;
mem[16'h72F3] = 8'h72;
mem[16'h72F4] = 8'hA9;
mem[16'h72F5] = 8'h12;
mem[16'h72F6] = 8'h8D;
mem[16'h72F7] = 8'h24;
mem[16'h72F8] = 8'h8C;
mem[16'h72F9] = 8'hA9;
mem[16'h72FA] = 8'h85;
mem[16'h72FB] = 8'hA0;
mem[16'h72FC] = 8'h4F;
mem[16'h72FD] = 8'h20;
mem[16'h72FE] = 8'h2B;
mem[16'h72FF] = 8'h8C;
mem[16'h7300] = 8'hBD;
mem[16'h7301] = 8'h2C;
mem[16'h7302] = 8'h5F;
mem[16'h7303] = 8'h85;
mem[16'h7304] = 8'h57;
mem[16'h7305] = 8'hBD;
mem[16'h7306] = 8'h1E;
mem[16'h7307] = 8'h5F;
mem[16'h7308] = 8'h85;
mem[16'h7309] = 8'h56;
mem[16'h730A] = 8'h20;
mem[16'h730B] = 8'hA8;
mem[16'h730C] = 8'h8B;
mem[16'h730D] = 8'h60;
mem[16'h730E] = 8'hA9;
mem[16'h730F] = 8'h26;
mem[16'h7310] = 8'hA0;
mem[16'h7311] = 8'h73;
mem[16'h7312] = 8'h20;
mem[16'h7313] = 8'h2B;
mem[16'h7314] = 8'h8C;
mem[16'h7315] = 8'hA9;
mem[16'h7316] = 8'h00;
mem[16'h7317] = 8'h85;
mem[16'h7318] = 8'h56;
mem[16'h7319] = 8'hA9;
mem[16'h731A] = 8'h78;
mem[16'h731B] = 8'h85;
mem[16'h731C] = 8'h57;
mem[16'h731D] = 8'hA9;
mem[16'h731E] = 8'h10;
mem[16'h731F] = 8'h8D;
mem[16'h7320] = 8'h24;
mem[16'h7321] = 8'h8C;
mem[16'h7322] = 8'h20;
mem[16'h7323] = 8'hA8;
mem[16'h7324] = 8'h8B;
mem[16'h7325] = 8'h60;
mem[16'h7326] = 8'h8C;
mem[16'h7327] = 8'h03;
mem[16'h7328] = 8'hDA;
mem[16'h7329] = 8'h05;
mem[16'h732A] = 8'hAA;
mem[16'h732B] = 8'h05;
mem[16'h732C] = 8'hAA;
mem[16'h732D] = 8'h05;
mem[16'h732E] = 8'hAC;
mem[16'h732F] = 8'h03;
mem[16'h7330] = 8'hA8;
mem[16'h7331] = 8'h02;
mem[16'h7332] = 8'hF0;
mem[16'h7333] = 8'h00;
mem[16'h7334] = 8'hA0;
mem[16'h7335] = 8'h00;
mem[16'h7336] = 8'hAE;
mem[16'h7337] = 8'h5A;
mem[16'h7338] = 8'h74;
mem[16'h7339] = 8'hCA;
mem[16'h733A] = 8'h30;
mem[16'h733B] = 8'h3B;
mem[16'h733C] = 8'h86;
mem[16'h733D] = 8'h70;
mem[16'h733E] = 8'hAD;
mem[16'h733F] = 8'h93;
mem[16'h7340] = 8'h73;
mem[16'h7341] = 8'hD0;
mem[16'h7342] = 8'h2F;
mem[16'h7343] = 8'h20;
mem[16'h7344] = 8'hA7;
mem[16'h7345] = 8'h73;
mem[16'h7346] = 8'hA6;
mem[16'h7347] = 8'h70;
mem[16'h7348] = 8'hBD;
mem[16'h7349] = 8'h84;
mem[16'h734A] = 8'h7B;
mem[16'h734B] = 8'h18;
mem[16'h734C] = 8'h69;
mem[16'h734D] = 8'h02;
mem[16'h734E] = 8'h9D;
mem[16'h734F] = 8'h84;
mem[16'h7350] = 8'h7B;
mem[16'h7351] = 8'hC9;
mem[16'h7352] = 8'hDB;
mem[16'h7353] = 8'h90;
mem[16'h7354] = 8'h23;
mem[16'h7355] = 8'h20;
mem[16'h7356] = 8'h8A;
mem[16'h7357] = 8'h7B;
mem[16'h7358] = 8'hAD;
mem[16'h7359] = 8'hB1;
mem[16'h735A] = 8'h4A;
mem[16'h735B] = 8'hF0;
mem[16'h735C] = 8'h06;
mem[16'h735D] = 8'hA9;
mem[16'h735E] = 8'h30;
mem[16'h735F] = 8'h8D;
mem[16'h7360] = 8'h93;
mem[16'h7361] = 8'h73;
mem[16'h7362] = 8'h60;
mem[16'h7363] = 8'hA6;
mem[16'h7364] = 8'h70;
mem[16'h7365] = 8'hA9;
mem[16'h7366] = 8'h01;
mem[16'h7367] = 8'h9D;
mem[16'h7368] = 8'h84;
mem[16'h7369] = 8'h7B;
mem[16'h736A] = 8'h20;
mem[16'h736B] = 8'h8A;
mem[16'h736C] = 8'h7B;
mem[16'h736D] = 8'hA6;
mem[16'h736E] = 8'h70;
mem[16'h736F] = 8'h4C;
mem[16'h7370] = 8'h78;
mem[16'h7371] = 8'h73;
mem[16'h7372] = 8'hCE;
mem[16'h7373] = 8'h93;
mem[16'h7374] = 8'h73;
mem[16'h7375] = 8'hF0;
mem[16'h7376] = 8'hEC;
mem[16'h7377] = 8'h60;
mem[16'h7378] = 8'hCE;
mem[16'h7379] = 8'h92;
mem[16'h737A] = 8'h73;
mem[16'h737B] = 8'hD0;
mem[16'h737C] = 8'hBC;
mem[16'h737D] = 8'hA9;
mem[16'h737E] = 8'h1E;
mem[16'h737F] = 8'h8D;
mem[16'h7380] = 8'h92;
mem[16'h7381] = 8'h73;
mem[16'h7382] = 8'h20;
mem[16'h7383] = 8'h94;
mem[16'h7384] = 8'h73;
mem[16'h7385] = 8'hAD;
mem[16'h7386] = 8'h0F;
mem[16'h7387] = 8'h7C;
mem[16'h7388] = 8'h49;
mem[16'h7389] = 8'h01;
mem[16'h738A] = 8'h8D;
mem[16'h738B] = 8'h0F;
mem[16'h738C] = 8'h7C;
mem[16'h738D] = 8'hA6;
mem[16'h738E] = 8'h70;
mem[16'h738F] = 8'h4C;
mem[16'h7390] = 8'h39;
mem[16'h7391] = 8'h73;
mem[16'h7392] = 8'h0F;
mem[16'h7393] = 8'h00;
mem[16'h7394] = 8'hAD;
mem[16'h7395] = 8'h0F;
mem[16'h7396] = 8'h7C;
mem[16'h7397] = 8'hD0;
mem[16'h7398] = 8'h07;
mem[16'h7399] = 8'h20;
mem[16'h739A] = 8'hED;
mem[16'h739B] = 8'h7B;
mem[16'h739C] = 8'h20;
mem[16'h739D] = 8'hCE;
mem[16'h739E] = 8'h7B;
mem[16'h739F] = 8'h60;
mem[16'h73A0] = 8'h20;
mem[16'h73A1] = 8'hCE;
mem[16'h73A2] = 8'h7B;
mem[16'h73A3] = 8'h20;
mem[16'h73A4] = 8'hED;
mem[16'h73A5] = 8'h7B;
mem[16'h73A6] = 8'h60;
mem[16'h73A7] = 8'hA6;
mem[16'h73A8] = 8'h70;
mem[16'h73A9] = 8'hBD;
mem[16'h73AA] = 8'h87;
mem[16'h73AB] = 8'h7B;
mem[16'h73AC] = 8'h18;
mem[16'h73AD] = 8'h69;
mem[16'h73AE] = 8'h04;
mem[16'h73AF] = 8'h85;
mem[16'h73B0] = 8'h56;
mem[16'h73B1] = 8'hBC;
mem[16'h73B2] = 8'h84;
mem[16'h73B3] = 8'h7B;
mem[16'h73B4] = 8'h84;
mem[16'h73B5] = 8'h57;
mem[16'h73B6] = 8'hB9;
mem[16'h73B7] = 8'h3E;
mem[16'h73B8] = 8'h8C;
mem[16'h73B9] = 8'hAA;
mem[16'h73BA] = 8'hBD;
mem[16'h73BB] = 8'h94;
mem[16'h73BC] = 8'h8E;
mem[16'h73BD] = 8'hAA;
mem[16'h73BE] = 8'hBD;
mem[16'h73BF] = 8'h5B;
mem[16'h73C0] = 8'h74;
mem[16'h73C1] = 8'hBC;
mem[16'h73C2] = 8'h62;
mem[16'h73C3] = 8'h74;
mem[16'h73C4] = 8'h20;
mem[16'h73C5] = 8'h0E;
mem[16'h73C6] = 8'h69;
mem[16'h73C7] = 8'hA9;
mem[16'h73C8] = 8'h1E;
mem[16'h73C9] = 8'h8D;
mem[16'h73CA] = 8'h07;
mem[16'h73CB] = 8'h69;
mem[16'h73CC] = 8'h20;
mem[16'h73CD] = 8'h9F;
mem[16'h73CE] = 8'h68;
mem[16'h73CF] = 8'hA6;
mem[16'h73D0] = 8'h70;
mem[16'h73D1] = 8'hBD;
mem[16'h73D2] = 8'h87;
mem[16'h73D3] = 8'h7B;
mem[16'h73D4] = 8'h18;
mem[16'h73D5] = 8'h69;
mem[16'h73D6] = 8'h02;
mem[16'h73D7] = 8'h85;
mem[16'h73D8] = 8'h56;
mem[16'h73D9] = 8'hBD;
mem[16'h73DA] = 8'h84;
mem[16'h73DB] = 8'h7B;
mem[16'h73DC] = 8'h18;
mem[16'h73DD] = 8'h69;
mem[16'h73DE] = 8'h15;
mem[16'h73DF] = 8'hA8;
mem[16'h73E0] = 8'h84;
mem[16'h73E1] = 8'h57;
mem[16'h73E2] = 8'hB9;
mem[16'h73E3] = 8'h3E;
mem[16'h73E4] = 8'h8C;
mem[16'h73E5] = 8'hAA;
mem[16'h73E6] = 8'hBD;
mem[16'h73E7] = 8'h94;
mem[16'h73E8] = 8'h8E;
mem[16'h73E9] = 8'hAA;
mem[16'h73EA] = 8'hBD;
mem[16'h73EB] = 8'h69;
mem[16'h73EC] = 8'h74;
mem[16'h73ED] = 8'hBC;
mem[16'h73EE] = 8'h70;
mem[16'h73EF] = 8'h74;
mem[16'h73F0] = 8'h20;
mem[16'h73F1] = 8'hD1;
mem[16'h73F2] = 8'h8A;
mem[16'h73F3] = 8'hA9;
mem[16'h73F4] = 8'h20;
mem[16'h73F5] = 8'h8D;
mem[16'h73F6] = 8'hCA;
mem[16'h73F7] = 8'h8A;
mem[16'h73F8] = 8'h20;
mem[16'h73F9] = 8'h79;
mem[16'h73FA] = 8'h8A;
mem[16'h73FB] = 8'hAD;
mem[16'h73FC] = 8'h0F;
mem[16'h73FD] = 8'h7C;
mem[16'h73FE] = 8'hD0;
mem[16'h73FF] = 8'h2D;
mem[16'h7400] = 8'hA6;
mem[16'h7401] = 8'h70;
mem[16'h7402] = 8'hBD;
mem[16'h7403] = 8'h87;
mem[16'h7404] = 8'h7B;
mem[16'h7405] = 8'h18;
mem[16'h7406] = 8'h69;
mem[16'h7407] = 8'h02;
mem[16'h7408] = 8'h85;
mem[16'h7409] = 8'h56;
mem[16'h740A] = 8'hBD;
mem[16'h740B] = 8'h84;
mem[16'h740C] = 8'h7B;
mem[16'h740D] = 8'h18;
mem[16'h740E] = 8'h69;
mem[16'h740F] = 8'h23;
mem[16'h7410] = 8'hA8;
mem[16'h7411] = 8'h84;
mem[16'h7412] = 8'h57;
mem[16'h7413] = 8'hB9;
mem[16'h7414] = 8'h3E;
mem[16'h7415] = 8'h8C;
mem[16'h7416] = 8'hAA;
mem[16'h7417] = 8'hBD;
mem[16'h7418] = 8'h94;
mem[16'h7419] = 8'h8E;
mem[16'h741A] = 8'hAA;
mem[16'h741B] = 8'hBD;
mem[16'h741C] = 8'h85;
mem[16'h741D] = 8'h74;
mem[16'h741E] = 8'hBC;
mem[16'h741F] = 8'h8C;
mem[16'h7420] = 8'h74;
mem[16'h7421] = 8'h20;
mem[16'h7422] = 8'hD1;
mem[16'h7423] = 8'h8A;
mem[16'h7424] = 8'hA9;
mem[16'h7425] = 8'h20;
mem[16'h7426] = 8'h8D;
mem[16'h7427] = 8'hCA;
mem[16'h7428] = 8'h8A;
mem[16'h7429] = 8'h20;
mem[16'h742A] = 8'h79;
mem[16'h742B] = 8'h8A;
mem[16'h742C] = 8'h60;
mem[16'h742D] = 8'hA6;
mem[16'h742E] = 8'h70;
mem[16'h742F] = 8'hBD;
mem[16'h7430] = 8'h87;
mem[16'h7431] = 8'h7B;
mem[16'h7432] = 8'h85;
mem[16'h7433] = 8'h56;
mem[16'h7434] = 8'hBD;
mem[16'h7435] = 8'h84;
mem[16'h7436] = 8'h7B;
mem[16'h7437] = 8'h18;
mem[16'h7438] = 8'h69;
mem[16'h7439] = 8'h23;
mem[16'h743A] = 8'hA8;
mem[16'h743B] = 8'h84;
mem[16'h743C] = 8'h57;
mem[16'h743D] = 8'hB9;
mem[16'h743E] = 8'h3E;
mem[16'h743F] = 8'h8C;
mem[16'h7440] = 8'hAA;
mem[16'h7441] = 8'hBD;
mem[16'h7442] = 8'h94;
mem[16'h7443] = 8'h8E;
mem[16'h7444] = 8'hAA;
mem[16'h7445] = 8'hBD;
mem[16'h7446] = 8'h77;
mem[16'h7447] = 8'h74;
mem[16'h7448] = 8'hBC;
mem[16'h7449] = 8'h7E;
mem[16'h744A] = 8'h74;
mem[16'h744B] = 8'h20;
mem[16'h744C] = 8'h3B;
mem[16'h744D] = 8'h8B;
mem[16'h744E] = 8'hA9;
mem[16'h744F] = 8'h1E;
mem[16'h7450] = 8'h8D;
mem[16'h7451] = 8'h34;
mem[16'h7452] = 8'h8B;
mem[16'h7453] = 8'h20;
mem[16'h7454] = 8'hF0;
mem[16'h7455] = 8'h8A;
mem[16'h7456] = 8'h60;
mem[16'h7457] = 8'hF0;
mem[16'h7458] = 8'hD4;
mem[16'h7459] = 8'h60;
mem[16'h745A] = 8'h00;
mem[16'h745B] = 8'h15;
mem[16'h745C] = 8'h33;
mem[16'h745D] = 8'h51;
mem[16'h745E] = 8'h6F;
mem[16'h745F] = 8'h8D;
mem[16'h7460] = 8'hAB;
mem[16'h7461] = 8'hC9;
mem[16'h7462] = 8'h87;
mem[16'h7463] = 8'h87;
mem[16'h7464] = 8'h87;
mem[16'h7465] = 8'h87;
mem[16'h7466] = 8'h87;
mem[16'h7467] = 8'h87;
mem[16'h7468] = 8'h87;
mem[16'h7469] = 8'hA7;
mem[16'h746A] = 8'h87;
mem[16'h746B] = 8'h67;
mem[16'h746C] = 8'h47;
mem[16'h746D] = 8'h27;
mem[16'h746E] = 8'h07;
mem[16'h746F] = 8'hE7;
mem[16'h7470] = 8'h88;
mem[16'h7471] = 8'h88;
mem[16'h7472] = 8'h88;
mem[16'h7473] = 8'h88;
mem[16'h7474] = 8'h88;
mem[16'h7475] = 8'h88;
mem[16'h7476] = 8'h87;
mem[16'h7477] = 8'h7B;
mem[16'h7478] = 8'h5D;
mem[16'h7479] = 8'h3F;
mem[16'h747A] = 8'h21;
mem[16'h747B] = 8'h03;
mem[16'h747C] = 8'hE5;
mem[16'h747D] = 8'hC7;
mem[16'h747E] = 8'h89;
mem[16'h747F] = 8'h89;
mem[16'h7480] = 8'h89;
mem[16'h7481] = 8'h89;
mem[16'h7482] = 8'h89;
mem[16'h7483] = 8'h88;
mem[16'h7484] = 8'h88;
mem[16'h7485] = 8'h59;
mem[16'h7486] = 8'h39;
mem[16'h7487] = 8'h19;
mem[16'h7488] = 8'hF9;
mem[16'h7489] = 8'hD9;
mem[16'h748A] = 8'hB9;
mem[16'h748B] = 8'h99;
mem[16'h748C] = 8'h8A;
mem[16'h748D] = 8'h8A;
mem[16'h748E] = 8'h8A;
mem[16'h748F] = 8'h89;
mem[16'h7490] = 8'h89;
mem[16'h7491] = 8'h89;
mem[16'h7492] = 8'h89;
mem[16'h7493] = 8'h5D;
mem[16'h7494] = 8'h01;
mem[16'h7495] = 8'h00;
mem[16'h7496] = 8'h00;
mem[16'h7497] = 8'h56;
mem[16'h7498] = 8'h03;
mem[16'h7499] = 8'h00;
mem[16'h749A] = 8'h00;
mem[16'h749B] = 8'h30;
mem[16'h749C] = 8'h03;
mem[16'h749D] = 8'h00;
mem[16'h749E] = 8'h00;
mem[16'h749F] = 8'h60;
mem[16'h74A0] = 8'h03;
mem[16'h74A1] = 8'h0F;
mem[16'h74A2] = 8'h00;
mem[16'h74A3] = 8'h40;
mem[16'h74A4] = 8'h47;
mem[16'h74A5] = 8'h19;
mem[16'h74A6] = 8'h00;
mem[16'h74A7] = 8'h00;
mem[16'h74A8] = 8'h6F;
mem[16'h74A9] = 8'h3F;
mem[16'h74AA] = 8'h00;
mem[16'h74AB] = 8'h00;
mem[16'h74AC] = 8'h46;
mem[16'h74AD] = 8'h79;
mem[16'h74AE] = 8'h00;
mem[16'h74AF] = 8'h00;
mem[16'h74B0] = 8'h6C;
mem[16'h74B1] = 8'h50;
mem[16'h74B2] = 8'h00;
mem[16'h74B3] = 8'h3A;
mem[16'h74B4] = 8'h03;
mem[16'h74B5] = 8'h00;
mem[16'h74B6] = 8'h00;
mem[16'h74B7] = 8'h2C;
mem[16'h74B8] = 8'h07;
mem[16'h74B9] = 8'h00;
mem[16'h74BA] = 8'h00;
mem[16'h74BB] = 8'h60;
mem[16'h74BC] = 8'h06;
mem[16'h74BD] = 8'h00;
mem[16'h74BE] = 8'h00;
mem[16'h74BF] = 8'h40;
mem[16'h74C0] = 8'h07;
mem[16'h74C1] = 8'h1E;
mem[16'h74C2] = 8'h00;
mem[16'h74C3] = 8'h00;
mem[16'h74C4] = 8'h0F;
mem[16'h74C5] = 8'h33;
mem[16'h74C6] = 8'h00;
mem[16'h74C7] = 8'h00;
mem[16'h74C8] = 8'h5E;
mem[16'h74C9] = 8'h7F;
mem[16'h74CA] = 8'h00;
mem[16'h74CB] = 8'h00;
mem[16'h74CC] = 8'h0C;
mem[16'h74CD] = 8'h73;
mem[16'h74CE] = 8'h01;
mem[16'h74CF] = 8'h00;
mem[16'h74D0] = 8'h58;
mem[16'h74D1] = 8'h21;
mem[16'h74D2] = 8'h01;
mem[16'h74D3] = 8'h74;
mem[16'h74D4] = 8'h06;
mem[16'h74D5] = 8'h00;
mem[16'h74D6] = 8'h00;
mem[16'h74D7] = 8'h58;
mem[16'h74D8] = 8'h0E;
mem[16'h74D9] = 8'h00;
mem[16'h74DA] = 8'h00;
mem[16'h74DB] = 8'h40;
mem[16'h74DC] = 8'h0D;
mem[16'h74DD] = 8'h00;
mem[16'h74DE] = 8'h00;
mem[16'h74DF] = 8'h00;
mem[16'h74E0] = 8'h0F;
mem[16'h74E1] = 8'h3C;
mem[16'h74E2] = 8'h00;
mem[16'h74E3] = 8'h00;
mem[16'h74E4] = 8'h1E;
mem[16'h74E5] = 8'h66;
mem[16'h74E6] = 8'h00;
mem[16'h74E7] = 8'h00;
mem[16'h74E8] = 8'h3C;
mem[16'h74E9] = 8'h7F;
mem[16'h74EA] = 8'h01;
mem[16'h74EB] = 8'h00;
mem[16'h74EC] = 8'h18;
mem[16'h74ED] = 8'h66;
mem[16'h74EE] = 8'h03;
mem[16'h74EF] = 8'h00;
mem[16'h74F0] = 8'h30;
mem[16'h74F1] = 8'h43;
mem[16'h74F2] = 8'h02;
mem[16'h74F3] = 8'h68;
mem[16'h74F4] = 8'h0D;
mem[16'h74F5] = 8'h00;
mem[16'h74F6] = 8'h00;
mem[16'h74F7] = 8'h30;
mem[16'h74F8] = 8'h1D;
mem[16'h74F9] = 8'h00;
mem[16'h74FA] = 8'h00;
mem[16'h74FB] = 8'h00;
mem[16'h74FC] = 8'h1B;
mem[16'h74FD] = 8'h00;
mem[16'h74FE] = 8'h00;
mem[16'h74FF] = 8'h00;
mem[16'h7500] = 8'h1E;
mem[16'h7501] = 8'h78;
mem[16'h7502] = 8'h00;
mem[16'h7503] = 8'h00;
mem[16'h7504] = 8'h3C;
mem[16'h7505] = 8'h4C;
mem[16'h7506] = 8'h01;
mem[16'h7507] = 8'h00;
mem[16'h7508] = 8'h78;
mem[16'h7509] = 8'h7E;
mem[16'h750A] = 8'h03;
mem[16'h750B] = 8'h00;
mem[16'h750C] = 8'h30;
mem[16'h750D] = 8'h4C;
mem[16'h750E] = 8'h07;
mem[16'h750F] = 8'h00;
mem[16'h7510] = 8'h60;
mem[16'h7511] = 8'h06;
mem[16'h7512] = 8'h05;
mem[16'h7513] = 8'h50;
mem[16'h7514] = 8'h1B;
mem[16'h7515] = 8'h00;
mem[16'h7516] = 8'h00;
mem[16'h7517] = 8'h60;
mem[16'h7518] = 8'h3A;
mem[16'h7519] = 8'h00;
mem[16'h751A] = 8'h00;
mem[16'h751B] = 8'h00;
mem[16'h751C] = 8'h36;
mem[16'h751D] = 8'h00;
mem[16'h751E] = 8'h00;
mem[16'h751F] = 8'h00;
mem[16'h7520] = 8'h3C;
mem[16'h7521] = 8'h70;
mem[16'h7522] = 8'h01;
mem[16'h7523] = 8'h00;
mem[16'h7524] = 8'h78;
mem[16'h7525] = 8'h18;
mem[16'h7526] = 8'h03;
mem[16'h7527] = 8'h00;
mem[16'h7528] = 8'h70;
mem[16'h7529] = 8'h7D;
mem[16'h752A] = 8'h07;
mem[16'h752B] = 8'h00;
mem[16'h752C] = 8'h60;
mem[16'h752D] = 8'h18;
mem[16'h752E] = 8'h0F;
mem[16'h752F] = 8'h00;
mem[16'h7530] = 8'h40;
mem[16'h7531] = 8'h0D;
mem[16'h7532] = 8'h0A;
mem[16'h7533] = 8'h20;
mem[16'h7534] = 8'h37;
mem[16'h7535] = 8'h00;
mem[16'h7536] = 8'h00;
mem[16'h7537] = 8'h40;
mem[16'h7538] = 8'h75;
mem[16'h7539] = 8'h00;
mem[16'h753A] = 8'h00;
mem[16'h753B] = 8'h00;
mem[16'h753C] = 8'h6C;
mem[16'h753D] = 8'h00;
mem[16'h753E] = 8'h00;
mem[16'h753F] = 8'h00;
mem[16'h7540] = 8'h78;
mem[16'h7541] = 8'h60;
mem[16'h7542] = 8'h03;
mem[16'h7543] = 8'h00;
mem[16'h7544] = 8'h70;
mem[16'h7545] = 8'h31;
mem[16'h7546] = 8'h06;
mem[16'h7547] = 8'h00;
mem[16'h7548] = 8'h60;
mem[16'h7549] = 8'h7B;
mem[16'h754A] = 8'h0F;
mem[16'h754B] = 8'h00;
mem[16'h754C] = 8'h40;
mem[16'h754D] = 8'h31;
mem[16'h754E] = 8'h1E;
mem[16'h754F] = 8'h00;
mem[16'h7550] = 8'h00;
mem[16'h7551] = 8'h1B;
mem[16'h7552] = 8'h14;
mem[16'h7553] = 8'h40;
mem[16'h7554] = 8'h6E;
mem[16'h7555] = 8'h00;
mem[16'h7556] = 8'h00;
mem[16'h7557] = 8'h00;
mem[16'h7558] = 8'h6B;
mem[16'h7559] = 8'h01;
mem[16'h755A] = 8'h00;
mem[16'h755B] = 8'h00;
mem[16'h755C] = 8'h58;
mem[16'h755D] = 8'h01;
mem[16'h755E] = 8'h00;
mem[16'h755F] = 8'h00;
mem[16'h7560] = 8'h70;
mem[16'h7561] = 8'h41;
mem[16'h7562] = 8'h07;
mem[16'h7563] = 8'h00;
mem[16'h7564] = 8'h60;
mem[16'h7565] = 8'h63;
mem[16'h7566] = 8'h0C;
mem[16'h7567] = 8'h00;
mem[16'h7568] = 8'h40;
mem[16'h7569] = 8'h77;
mem[16'h756A] = 8'h1F;
mem[16'h756B] = 8'h00;
mem[16'h756C] = 8'h00;
mem[16'h756D] = 8'h63;
mem[16'h756E] = 8'h3C;
mem[16'h756F] = 8'h00;
mem[16'h7570] = 8'h00;
mem[16'h7571] = 8'h36;
mem[16'h7572] = 8'h28;
mem[16'h7573] = 8'h00;
mem[16'h7574] = 8'h04;
mem[16'h7575] = 8'h28;
mem[16'h7576] = 8'h40;
mem[16'h7577] = 8'h60;
mem[16'h7578] = 8'h17;
mem[16'h7579] = 8'h1E;
mem[16'h757A] = 8'h58;
mem[16'h757B] = 8'h17;
mem[16'h757C] = 8'h30;
mem[16'h757D] = 8'h17;
mem[16'h757E] = 8'h30;
mem[16'h757F] = 8'h17;
mem[16'h7580] = 8'h30;
mem[16'h7581] = 8'h1E;
mem[16'h7582] = 8'h58;
mem[16'h7583] = 8'h60;
mem[16'h7584] = 8'h17;
mem[16'h7585] = 8'h28;
mem[16'h7586] = 8'h40;
mem[16'h7587] = 8'h00;
mem[16'h7588] = 8'h04;
mem[16'h7589] = 8'h20;
mem[16'h758A] = 8'h05;
mem[16'h758B] = 8'h08;
mem[16'h758C] = 8'h10;
mem[16'h758D] = 8'h20;
mem[16'h758E] = 8'h05;
mem[16'h758F] = 8'h62;
mem[16'h7590] = 8'h47;
mem[16'h7591] = 8'h3A;
mem[16'h7592] = 8'h5C;
mem[16'h7593] = 8'h1A;
mem[16'h7594] = 8'h58;
mem[16'h7595] = 8'h3A;
mem[16'h7596] = 8'h5C;
mem[16'h7597] = 8'h62;
mem[16'h7598] = 8'h47;
mem[16'h7599] = 8'h20;
mem[16'h759A] = 8'h05;
mem[16'h759B] = 8'h08;
mem[16'h759C] = 8'h10;
mem[16'h759D] = 8'h20;
mem[16'h759E] = 8'h05;
mem[16'h759F] = 8'h00;
mem[16'h75A0] = 8'h00;
mem[16'h75A1] = 8'h00;
mem[16'h75A2] = 8'h00;
mem[16'h75A3] = 8'h20;
mem[16'h75A4] = 8'h05;
mem[16'h75A5] = 8'h00;
mem[16'h75A6] = 8'h00;
mem[16'h75A7] = 8'h48;
mem[16'h75A8] = 8'h13;
mem[16'h75A9] = 8'h68;
mem[16'h75AA] = 8'h17;
mem[16'h75AB] = 8'h48;
mem[16'h75AC] = 8'h13;
mem[16'h75AD] = 8'h00;
mem[16'h75AE] = 8'h00;
mem[16'h75AF] = 8'h20;
mem[16'h75B0] = 8'h05;
mem[16'h75B1] = 8'hA9;
mem[16'h75B2] = 8'h73;
mem[16'h75B3] = 8'hA0;
mem[16'h75B4] = 8'h75;
mem[16'h75B5] = 8'h20;
mem[16'h75B6] = 8'h2B;
mem[16'h75B7] = 8'h8C;
mem[16'h75B8] = 8'hA9;
mem[16'h75B9] = 8'h16;
mem[16'h75BA] = 8'h8D;
mem[16'h75BB] = 8'h24;
mem[16'h75BC] = 8'h8C;
mem[16'h75BD] = 8'hA6;
mem[16'h75BE] = 8'h70;
mem[16'h75BF] = 8'hBD;
mem[16'h75C0] = 8'h2C;
mem[16'h75C1] = 8'h5F;
mem[16'h75C2] = 8'h85;
mem[16'h75C3] = 8'h57;
mem[16'h75C4] = 8'hBD;
mem[16'h75C5] = 8'h1E;
mem[16'h75C6] = 8'h5F;
mem[16'h75C7] = 8'h85;
mem[16'h75C8] = 8'h56;
mem[16'h75C9] = 8'h20;
mem[16'h75CA] = 8'hA8;
mem[16'h75CB] = 8'h8B;
mem[16'h75CC] = 8'h60;
mem[16'h75CD] = 8'hA9;
mem[16'h75CE] = 8'h89;
mem[16'h75CF] = 8'hA0;
mem[16'h75D0] = 8'h75;
mem[16'h75D1] = 8'h20;
mem[16'h75D2] = 8'h2B;
mem[16'h75D3] = 8'h8C;
mem[16'h75D4] = 8'hA9;
mem[16'h75D5] = 8'h16;
mem[16'h75D6] = 8'h8D;
mem[16'h75D7] = 8'h24;
mem[16'h75D8] = 8'h8C;
mem[16'h75D9] = 8'h4C;
mem[16'h75DA] = 8'hBD;
mem[16'h75DB] = 8'h75;
mem[16'h75DC] = 8'hA9;
mem[16'h75DD] = 8'h9F;
mem[16'h75DE] = 8'hA0;
mem[16'h75DF] = 8'h75;
mem[16'h75E0] = 8'h20;
mem[16'h75E1] = 8'h2B;
mem[16'h75E2] = 8'h8C;
mem[16'h75E3] = 8'hA9;
mem[16'h75E4] = 8'h12;
mem[16'h75E5] = 8'h8D;
mem[16'h75E6] = 8'h24;
mem[16'h75E7] = 8'h8C;
mem[16'h75E8] = 8'h4C;
mem[16'h75E9] = 8'hBD;
mem[16'h75EA] = 8'h75;
mem[16'h75EB] = 8'hA6;
mem[16'h75EC] = 8'h70;
mem[16'h75ED] = 8'hBD;
mem[16'h75EE] = 8'h1E;
mem[16'h75EF] = 8'h5F;
mem[16'h75F0] = 8'h85;
mem[16'h75F1] = 8'h56;
mem[16'h75F2] = 8'hBC;
mem[16'h75F3] = 8'h2C;
mem[16'h75F4] = 8'h5F;
mem[16'h75F5] = 8'h84;
mem[16'h75F6] = 8'h57;
mem[16'h75F7] = 8'hB9;
mem[16'h75F8] = 8'h3E;
mem[16'h75F9] = 8'h8C;
mem[16'h75FA] = 8'hAA;
mem[16'h75FB] = 8'hBD;
mem[16'h75FC] = 8'h94;
mem[16'h75FD] = 8'h8E;
mem[16'h75FE] = 8'hAA;
mem[16'h75FF] = 8'hBD;
mem[16'h7600] = 8'h37;
mem[16'h7601] = 8'h76;
mem[16'h7602] = 8'hBC;
mem[16'h7603] = 8'h3E;
mem[16'h7604] = 8'h76;
mem[16'h7605] = 8'h20;
mem[16'h7606] = 8'hD1;
mem[16'h7607] = 8'h8A;
mem[16'h7608] = 8'hA9;
mem[16'h7609] = 8'h2C;
mem[16'h760A] = 8'h8D;
mem[16'h760B] = 8'hCA;
mem[16'h760C] = 8'h8A;
mem[16'h760D] = 8'h20;
mem[16'h760E] = 8'h79;
mem[16'h760F] = 8'h8A;
mem[16'h7610] = 8'h60;
mem[16'h7611] = 8'hA6;
mem[16'h7612] = 8'h70;
mem[16'h7613] = 8'hBD;
mem[16'h7614] = 8'h1E;
mem[16'h7615] = 8'h5F;
mem[16'h7616] = 8'h85;
mem[16'h7617] = 8'h56;
mem[16'h7618] = 8'hBC;
mem[16'h7619] = 8'h2C;
mem[16'h761A] = 8'h5F;
mem[16'h761B] = 8'h84;
mem[16'h761C] = 8'h57;
mem[16'h761D] = 8'hB9;
mem[16'h761E] = 8'h3E;
mem[16'h761F] = 8'h8C;
mem[16'h7620] = 8'hAA;
mem[16'h7621] = 8'hBD;
mem[16'h7622] = 8'h94;
mem[16'h7623] = 8'h8E;
mem[16'h7624] = 8'hAA;
mem[16'h7625] = 8'hBD;
mem[16'h7626] = 8'h45;
mem[16'h7627] = 8'h76;
mem[16'h7628] = 8'hBC;
mem[16'h7629] = 8'h4C;
mem[16'h762A] = 8'h76;
mem[16'h762B] = 8'h20;
mem[16'h762C] = 8'hD1;
mem[16'h762D] = 8'h8A;
mem[16'h762E] = 8'hA9;
mem[16'h762F] = 8'h24;
mem[16'h7630] = 8'h8D;
mem[16'h7631] = 8'hCA;
mem[16'h7632] = 8'h8A;
mem[16'h7633] = 8'h20;
mem[16'h7634] = 8'h79;
mem[16'h7635] = 8'h8A;
mem[16'h7636] = 8'h60;
mem[16'h7637] = 8'h6E;
mem[16'h7638] = 8'h9A;
mem[16'h7639] = 8'hC6;
mem[16'h763A] = 8'hF2;
mem[16'h763B] = 8'h1E;
mem[16'h763C] = 8'h4A;
mem[16'h763D] = 8'h76;
mem[16'h763E] = 8'h81;
mem[16'h763F] = 8'h81;
mem[16'h7640] = 8'h81;
mem[16'h7641] = 8'h81;
mem[16'h7642] = 8'h82;
mem[16'h7643] = 8'h82;
mem[16'h7644] = 8'h82;
mem[16'h7645] = 8'h3B;
mem[16'h7646] = 8'h5F;
mem[16'h7647] = 8'h83;
mem[16'h7648] = 8'hA7;
mem[16'h7649] = 8'hCB;
mem[16'h764A] = 8'hEF;
mem[16'h764B] = 8'h13;
mem[16'h764C] = 8'h84;
mem[16'h764D] = 8'h84;
mem[16'h764E] = 8'h84;
mem[16'h764F] = 8'h84;
mem[16'h7650] = 8'h84;
mem[16'h7651] = 8'h84;
mem[16'h7652] = 8'h85;
mem[16'h7653] = 8'h00;
mem[16'h7654] = 8'h00;
mem[16'h7655] = 8'h00;
mem[16'h7656] = 8'h00;
mem[16'h7657] = 8'h00;
mem[16'h7658] = 8'h00;
mem[16'h7659] = 8'h00;
mem[16'h765A] = 8'h00;
mem[16'h765B] = 8'h00;
mem[16'h765C] = 8'h00;
mem[16'h765D] = 8'h00;
mem[16'h765E] = 8'h00;
mem[16'h765F] = 8'h00;
mem[16'h7660] = 8'h00;
mem[16'h7661] = 8'h00;
mem[16'h7662] = 8'h00;
mem[16'h7663] = 8'h00;
mem[16'h7664] = 8'h00;
mem[16'h7665] = 8'h00;
mem[16'h7666] = 8'h0C;
mem[16'h7667] = 8'h00;
mem[16'h7668] = 8'h00;
mem[16'h7669] = 8'h12;
mem[16'h766A] = 8'h00;
mem[16'h766B] = 8'h00;
mem[16'h766C] = 8'h21;
mem[16'h766D] = 8'h00;
mem[16'h766E] = 8'h00;
mem[16'h766F] = 8'h21;
mem[16'h7670] = 8'h00;
mem[16'h7671] = 8'h00;
mem[16'h7672] = 8'h12;
mem[16'h7673] = 8'h00;
mem[16'h7674] = 8'h00;
mem[16'h7675] = 8'h0C;
mem[16'h7676] = 8'h00;
mem[16'h7677] = 8'h00;
mem[16'h7678] = 8'h00;
mem[16'h7679] = 8'h00;
mem[16'h767A] = 8'h00;
mem[16'h767B] = 8'h00;
mem[16'h767C] = 8'h00;
mem[16'h767D] = 8'h00;
mem[16'h767E] = 8'h00;
mem[16'h767F] = 8'h00;
mem[16'h7680] = 8'h00;
mem[16'h7681] = 8'h00;
mem[16'h7682] = 8'h00;
mem[16'h7683] = 8'h00;
mem[16'h7684] = 8'h00;
mem[16'h7685] = 8'h00;
mem[16'h7686] = 8'h00;
mem[16'h7687] = 8'h00;
mem[16'h7688] = 8'h00;
mem[16'h7689] = 8'h00;
mem[16'h768A] = 8'h00;
mem[16'h768B] = 8'h00;
mem[16'h768C] = 8'h00;
mem[16'h768D] = 8'h00;
mem[16'h768E] = 8'h00;
mem[16'h768F] = 8'h00;
mem[16'h7690] = 8'h00;
mem[16'h7691] = 8'h00;
mem[16'h7692] = 8'h00;
mem[16'h7693] = 8'h00;
mem[16'h7694] = 8'h00;
mem[16'h7695] = 8'h00;
mem[16'h7696] = 8'h1E;
mem[16'h7697] = 8'h00;
mem[16'h7698] = 8'h00;
mem[16'h7699] = 8'h21;
mem[16'h769A] = 8'h00;
mem[16'h769B] = 8'h40;
mem[16'h769C] = 8'h4C;
mem[16'h769D] = 8'h00;
mem[16'h769E] = 8'h20;
mem[16'h769F] = 8'h12;
mem[16'h76A0] = 8'h01;
mem[16'h76A1] = 8'h20;
mem[16'h76A2] = 8'h21;
mem[16'h76A3] = 8'h01;
mem[16'h76A4] = 8'h20;
mem[16'h76A5] = 8'h21;
mem[16'h76A6] = 8'h01;
mem[16'h76A7] = 8'h20;
mem[16'h76A8] = 8'h12;
mem[16'h76A9] = 8'h01;
mem[16'h76AA] = 8'h40;
mem[16'h76AB] = 8'h4C;
mem[16'h76AC] = 8'h00;
mem[16'h76AD] = 8'h00;
mem[16'h76AE] = 8'h21;
mem[16'h76AF] = 8'h00;
mem[16'h76B0] = 8'h00;
mem[16'h76B1] = 8'h1E;
mem[16'h76B2] = 8'h00;
mem[16'h76B3] = 8'h00;
mem[16'h76B4] = 8'h00;
mem[16'h76B5] = 8'h00;
mem[16'h76B6] = 8'h00;
mem[16'h76B7] = 8'h00;
mem[16'h76B8] = 8'h00;
mem[16'h76B9] = 8'h00;
mem[16'h76BA] = 8'h00;
mem[16'h76BB] = 8'h00;
mem[16'h76BC] = 8'h00;
mem[16'h76BD] = 8'h00;
mem[16'h76BE] = 8'h00;
mem[16'h76BF] = 8'h00;
mem[16'h76C0] = 8'h00;
mem[16'h76C1] = 8'h00;
mem[16'h76C2] = 8'h00;
mem[16'h76C3] = 8'h00;
mem[16'h76C4] = 8'h00;
mem[16'h76C5] = 8'h00;
mem[16'h76C6] = 8'h3F;
mem[16'h76C7] = 8'h00;
mem[16'h76C8] = 8'h40;
mem[16'h76C9] = 8'h40;
mem[16'h76CA] = 8'h00;
mem[16'h76CB] = 8'h20;
mem[16'h76CC] = 8'h1E;
mem[16'h76CD] = 8'h01;
mem[16'h76CE] = 8'h10;
mem[16'h76CF] = 8'h21;
mem[16'h76D0] = 8'h02;
mem[16'h76D1] = 8'h48;
mem[16'h76D2] = 8'h40;
mem[16'h76D3] = 8'h04;
mem[16'h76D4] = 8'h28;
mem[16'h76D5] = 8'h00;
mem[16'h76D6] = 8'h05;
mem[16'h76D7] = 8'h28;
mem[16'h76D8] = 8'h00;
mem[16'h76D9] = 8'h05;
mem[16'h76DA] = 8'h28;
mem[16'h76DB] = 8'h00;
mem[16'h76DC] = 8'h05;
mem[16'h76DD] = 8'h28;
mem[16'h76DE] = 8'h00;
mem[16'h76DF] = 8'h05;
mem[16'h76E0] = 8'h48;
mem[16'h76E1] = 8'h40;
mem[16'h76E2] = 8'h04;
mem[16'h76E3] = 8'h10;
mem[16'h76E4] = 8'h21;
mem[16'h76E5] = 8'h02;
mem[16'h76E6] = 8'h20;
mem[16'h76E7] = 8'h1E;
mem[16'h76E8] = 8'h01;
mem[16'h76E9] = 8'h40;
mem[16'h76EA] = 8'h40;
mem[16'h76EB] = 8'h00;
mem[16'h76EC] = 8'h00;
mem[16'h76ED] = 8'h3F;
mem[16'h76EE] = 8'h00;
mem[16'h76EF] = 8'h00;
mem[16'h76F0] = 8'h00;
mem[16'h76F1] = 8'h00;
mem[16'h76F2] = 8'h00;
mem[16'h76F3] = 8'h00;
mem[16'h76F4] = 8'h00;
mem[16'h76F5] = 8'h40;
mem[16'h76F6] = 8'h7F;
mem[16'h76F7] = 8'h00;
mem[16'h76F8] = 8'h20;
mem[16'h76F9] = 8'h00;
mem[16'h76FA] = 8'h01;
mem[16'h76FB] = 8'h10;
mem[16'h76FC] = 8'h3F;
mem[16'h76FD] = 8'h02;
mem[16'h76FE] = 8'h48;
mem[16'h76FF] = 8'h40;
mem[16'h7700] = 8'h04;
mem[16'h7701] = 8'h24;
mem[16'h7702] = 8'h00;
mem[16'h7703] = 8'h09;
mem[16'h7704] = 8'h12;
mem[16'h7705] = 8'h00;
mem[16'h7706] = 8'h12;
mem[16'h7707] = 8'h0A;
mem[16'h7708] = 8'h00;
mem[16'h7709] = 8'h14;
mem[16'h770A] = 8'h0A;
mem[16'h770B] = 8'h00;
mem[16'h770C] = 8'h14;
mem[16'h770D] = 8'h0A;
mem[16'h770E] = 8'h00;
mem[16'h770F] = 8'h14;
mem[16'h7710] = 8'h0A;
mem[16'h7711] = 8'h00;
mem[16'h7712] = 8'h14;
mem[16'h7713] = 8'h0A;
mem[16'h7714] = 8'h00;
mem[16'h7715] = 8'h14;
mem[16'h7716] = 8'h0A;
mem[16'h7717] = 8'h00;
mem[16'h7718] = 8'h14;
mem[16'h7719] = 8'h12;
mem[16'h771A] = 8'h00;
mem[16'h771B] = 8'h12;
mem[16'h771C] = 8'h24;
mem[16'h771D] = 8'h00;
mem[16'h771E] = 8'h09;
mem[16'h771F] = 8'h48;
mem[16'h7720] = 8'h40;
mem[16'h7721] = 8'h04;
mem[16'h7722] = 8'h10;
mem[16'h7723] = 8'h3F;
mem[16'h7724] = 8'h02;
mem[16'h7725] = 8'h20;
mem[16'h7726] = 8'h00;
mem[16'h7727] = 8'h01;
mem[16'h7728] = 8'h40;
mem[16'h7729] = 8'h7F;
mem[16'h772A] = 8'h00;
mem[16'h772B] = 8'h40;
mem[16'h772C] = 8'h7F;
mem[16'h772D] = 8'h00;
mem[16'h772E] = 8'h20;
mem[16'h772F] = 8'h00;
mem[16'h7730] = 8'h01;
mem[16'h7731] = 8'h10;
mem[16'h7732] = 8'h00;
mem[16'h7733] = 8'h02;
mem[16'h7734] = 8'h08;
mem[16'h7735] = 8'h00;
mem[16'h7736] = 8'h04;
mem[16'h7737] = 8'h04;
mem[16'h7738] = 8'h00;
mem[16'h7739] = 8'h08;
mem[16'h773A] = 8'h02;
mem[16'h773B] = 8'h00;
mem[16'h773C] = 8'h10;
mem[16'h773D] = 8'h02;
mem[16'h773E] = 8'h00;
mem[16'h773F] = 8'h10;
mem[16'h7740] = 8'h02;
mem[16'h7741] = 8'h00;
mem[16'h7742] = 8'h10;
mem[16'h7743] = 8'h02;
mem[16'h7744] = 8'h00;
mem[16'h7745] = 8'h10;
mem[16'h7746] = 8'h02;
mem[16'h7747] = 8'h00;
mem[16'h7748] = 8'h10;
mem[16'h7749] = 8'h02;
mem[16'h774A] = 8'h00;
mem[16'h774B] = 8'h10;
mem[16'h774C] = 8'h02;
mem[16'h774D] = 8'h00;
mem[16'h774E] = 8'h10;
mem[16'h774F] = 8'h02;
mem[16'h7750] = 8'h00;
mem[16'h7751] = 8'h10;
mem[16'h7752] = 8'h04;
mem[16'h7753] = 8'h00;
mem[16'h7754] = 8'h08;
mem[16'h7755] = 8'h08;
mem[16'h7756] = 8'h00;
mem[16'h7757] = 8'h04;
mem[16'h7758] = 8'h10;
mem[16'h7759] = 8'h00;
mem[16'h775A] = 8'h02;
mem[16'h775B] = 8'h20;
mem[16'h775C] = 8'h00;
mem[16'h775D] = 8'h01;
mem[16'h775E] = 8'h40;
mem[16'h775F] = 8'h7F;
mem[16'h7760] = 8'h00;
mem[16'h7761] = 8'hAD;
mem[16'h7762] = 8'hC0;
mem[16'h7763] = 8'h62;
mem[16'h7764] = 8'h18;
mem[16'h7765] = 8'h6D;
mem[16'h7766] = 8'hC2;
mem[16'h7767] = 8'h62;
mem[16'h7768] = 8'h6D;
mem[16'h7769] = 8'hC1;
mem[16'h776A] = 8'h62;
mem[16'h776B] = 8'h6D;
mem[16'h776C] = 8'hC3;
mem[16'h776D] = 8'h62;
mem[16'h776E] = 8'hCD;
mem[16'h776F] = 8'hC7;
mem[16'h7770] = 8'h77;
mem[16'h7771] = 8'hB0;
mem[16'h7772] = 8'h14;
mem[16'h7773] = 8'hAD;
mem[16'h7774] = 8'h13;
mem[16'h7775] = 8'h87;
mem[16'h7776] = 8'h29;
mem[16'h7777] = 8'h0F;
mem[16'h7778] = 8'hC9;
mem[16'h7779] = 8'h08;
mem[16'h777A] = 8'h90;
mem[16'h777B] = 8'h0C;
mem[16'h777C] = 8'h29;
mem[16'h777D] = 8'h07;
mem[16'h777E] = 8'hAA;
mem[16'h777F] = 8'hAD;
mem[16'h7780] = 8'hC2;
mem[16'h7781] = 8'h62;
mem[16'h7782] = 8'hD0;
mem[16'h7783] = 8'h03;
mem[16'h7784] = 8'h20;
mem[16'h7785] = 8'h82;
mem[16'h7786] = 8'h62;
mem[16'h7787] = 8'h60;
mem[16'h7788] = 8'hAA;
mem[16'h7789] = 8'hAD;
mem[16'h778A] = 8'hC0;
mem[16'h778B] = 8'h62;
mem[16'h778C] = 8'hD0;
mem[16'h778D] = 8'hF9;
mem[16'h778E] = 8'hBD;
mem[16'h778F] = 8'hC8;
mem[16'h7790] = 8'h77;
mem[16'h7791] = 8'hC9;
mem[16'h7792] = 8'h33;
mem[16'h7793] = 8'hD0;
mem[16'h7794] = 8'h15;
mem[16'h7795] = 8'h8D;
mem[16'h7796] = 8'hBA;
mem[16'h7797] = 8'h62;
mem[16'h7798] = 8'hA9;
mem[16'h7799] = 8'h01;
mem[16'h779A] = 8'h8D;
mem[16'h779B] = 8'hD9;
mem[16'h779C] = 8'h77;
mem[16'h779D] = 8'hAD;
mem[16'h779E] = 8'h10;
mem[16'h779F] = 8'h51;
mem[16'h77A0] = 8'h38;
mem[16'h77A1] = 8'hED;
mem[16'h77A2] = 8'h16;
mem[16'h77A3] = 8'h51;
mem[16'h77A4] = 8'h8D;
mem[16'h77A5] = 8'hB8;
mem[16'h77A6] = 8'h62;
mem[16'h77A7] = 8'h4C;
mem[16'h77A8] = 8'hB6;
mem[16'h77A9] = 8'h77;
mem[16'h77AA] = 8'h8D;
mem[16'h77AB] = 8'hBA;
mem[16'h77AC] = 8'h62;
mem[16'h77AD] = 8'h8D;
mem[16'h77AE] = 8'hD8;
mem[16'h77AF] = 8'h77;
mem[16'h77B0] = 8'hBD;
mem[16'h77B1] = 8'hD0;
mem[16'h77B2] = 8'h77;
mem[16'h77B3] = 8'h8D;
mem[16'h77B4] = 8'hB8;
mem[16'h77B5] = 8'h62;
mem[16'h77B6] = 8'hA9;
mem[16'h77B7] = 8'h01;
mem[16'h77B8] = 8'h8D;
mem[16'h77B9] = 8'hC0;
mem[16'h77BA] = 8'h62;
mem[16'h77BB] = 8'hEE;
mem[16'h77BC] = 8'hC6;
mem[16'h77BD] = 8'h77;
mem[16'h77BE] = 8'hA9;
mem[16'h77BF] = 8'h00;
mem[16'h77C0] = 8'h85;
mem[16'h77C1] = 8'h70;
mem[16'h77C2] = 8'h20;
mem[16'h77C3] = 8'hF8;
mem[16'h77C4] = 8'h62;
mem[16'h77C5] = 8'h60;
mem[16'h77C6] = 8'h00;
mem[16'h77C7] = 8'h00;
mem[16'h77C8] = 8'h33;
mem[16'h77C9] = 8'h5E;
mem[16'h77CA] = 8'h5E;
mem[16'h77CB] = 8'h5E;
mem[16'h77CC] = 8'h5E;
mem[16'h77CD] = 8'h5E;
mem[16'h77CE] = 8'h33;
mem[16'h77CF] = 8'h5E;
mem[16'h77D0] = 8'h00;
mem[16'h77D1] = 8'h00;
mem[16'h77D2] = 8'h04;
mem[16'h77D3] = 8'h00;
mem[16'h77D4] = 8'h0C;
mem[16'h77D5] = 8'h1E;
mem[16'h77D6] = 8'h10;
mem[16'h77D7] = 8'h18;
mem[16'h77D8] = 8'h00;
mem[16'h77D9] = 8'h00;
mem[16'h77DA] = 8'hAD;
mem[16'h77DB] = 8'h33;
mem[16'h77DC] = 8'h7B;
mem[16'h77DD] = 8'hF0;
mem[16'h77DE] = 8'h0C;
mem[16'h77DF] = 8'h20;
mem[16'h77E0] = 8'hF4;
mem[16'h77E1] = 8'h77;
mem[16'h77E2] = 8'hAD;
mem[16'h77E3] = 8'h63;
mem[16'h77E4] = 8'h79;
mem[16'h77E5] = 8'hCD;
mem[16'h77E6] = 8'h13;
mem[16'h77E7] = 8'h51;
mem[16'h77E8] = 8'hF0;
mem[16'h77E9] = 8'h01;
mem[16'h77EA] = 8'h60;
mem[16'h77EB] = 8'hAD;
mem[16'h77EC] = 8'h33;
mem[16'h77ED] = 8'h7B;
mem[16'h77EE] = 8'hF0;
mem[16'h77EF] = 8'h03;
mem[16'h77F0] = 8'h20;
mem[16'h77F1] = 8'hF4;
mem[16'h77F2] = 8'h77;
mem[16'h77F3] = 8'h60;
mem[16'h77F4] = 8'hAD;
mem[16'h77F5] = 8'h63;
mem[16'h77F6] = 8'h79;
mem[16'h77F7] = 8'hCD;
mem[16'h77F8] = 8'h1E;
mem[16'h77F9] = 8'h5F;
mem[16'h77FA] = 8'hD0;
mem[16'h77FB] = 8'h03;
mem[16'h77FC] = 8'h4C;
mem[16'h77FD] = 8'h8E;
mem[16'h77FE] = 8'h78;
mem[16'h77FF] = 8'hCD;
mem[16'h7800] = 8'h26;
mem[16'h7801] = 8'h5F;
mem[16'h7802] = 8'hD0;
mem[16'h7803] = 8'h03;
mem[16'h7804] = 8'h4C;
mem[16'h7805] = 8'h8E;
mem[16'h7806] = 8'h78;
mem[16'h7807] = 8'h20;
mem[16'h7808] = 8'hE4;
mem[16'h7809] = 8'h78;
mem[16'h780A] = 8'hAE;
mem[16'h780B] = 8'h34;
mem[16'h780C] = 8'h7B;
mem[16'h780D] = 8'hAD;
mem[16'h780E] = 8'h63;
mem[16'h780F] = 8'h79;
mem[16'h7810] = 8'hCD;
mem[16'h7811] = 8'h03;
mem[16'h7812] = 8'h54;
mem[16'h7813] = 8'hD0;
mem[16'h7814] = 8'h0C;
mem[16'h7815] = 8'hBD;
mem[16'h7816] = 8'h00;
mem[16'h7817] = 8'h54;
mem[16'h7818] = 8'hFD;
mem[16'h7819] = 8'h0D;
mem[16'h781A] = 8'h54;
mem[16'h781B] = 8'h8D;
mem[16'h781C] = 8'hE3;
mem[16'h781D] = 8'h78;
mem[16'h781E] = 8'h4C;
mem[16'h781F] = 8'h3B;
mem[16'h7820] = 8'h78;
mem[16'h7821] = 8'hCD;
mem[16'h7822] = 8'h13;
mem[16'h7823] = 8'h51;
mem[16'h7824] = 8'hD0;
mem[16'h7825] = 8'h0C;
mem[16'h7826] = 8'hBD;
mem[16'h7827] = 8'h10;
mem[16'h7828] = 8'h51;
mem[16'h7829] = 8'hFD;
mem[16'h782A] = 8'h16;
mem[16'h782B] = 8'h51;
mem[16'h782C] = 8'h8D;
mem[16'h782D] = 8'hE3;
mem[16'h782E] = 8'h78;
mem[16'h782F] = 8'h4C;
mem[16'h7830] = 8'h3B;
mem[16'h7831] = 8'h78;
mem[16'h7832] = 8'hBD;
mem[16'h7833] = 8'h1F;
mem[16'h7834] = 8'h53;
mem[16'h7835] = 8'hFD;
mem[16'h7836] = 8'h28;
mem[16'h7837] = 8'h53;
mem[16'h7838] = 8'h8D;
mem[16'h7839] = 8'hE3;
mem[16'h783A] = 8'h78;
mem[16'h783B] = 8'hAD;
mem[16'h783C] = 8'h62;
mem[16'h783D] = 8'h79;
mem[16'h783E] = 8'h18;
mem[16'h783F] = 8'h69;
mem[16'h7840] = 8'h02;
mem[16'h7841] = 8'h8D;
mem[16'h7842] = 8'h62;
mem[16'h7843] = 8'h79;
mem[16'h7844] = 8'h69;
mem[16'h7845] = 8'h0B;
mem[16'h7846] = 8'hCD;
mem[16'h7847] = 8'hE3;
mem[16'h7848] = 8'h78;
mem[16'h7849] = 8'hB0;
mem[16'h784A] = 8'h13;
mem[16'h784B] = 8'hC9;
mem[16'h784C] = 8'hFC;
mem[16'h784D] = 8'h90;
mem[16'h784E] = 8'h0E;
mem[16'h784F] = 8'h20;
mem[16'h7850] = 8'h48;
mem[16'h7851] = 8'h79;
mem[16'h7852] = 8'hA9;
mem[16'h7853] = 8'h00;
mem[16'h7854] = 8'h8D;
mem[16'h7855] = 8'h33;
mem[16'h7856] = 8'h7B;
mem[16'h7857] = 8'hAD;
mem[16'h7858] = 8'hDF;
mem[16'h7859] = 8'h91;
mem[16'h785A] = 8'h8D;
mem[16'h785B] = 8'hDB;
mem[16'h785C] = 8'h91;
mem[16'h785D] = 8'h60;
mem[16'h785E] = 8'h38;
mem[16'h785F] = 8'hED;
mem[16'h7860] = 8'hCF;
mem[16'h7861] = 8'h4D;
mem[16'h7862] = 8'h20;
mem[16'h7863] = 8'h62;
mem[16'h7864] = 8'h65;
mem[16'h7865] = 8'hC9;
mem[16'h7866] = 8'h04;
mem[16'h7867] = 8'hB0;
mem[16'h7868] = 8'h16;
mem[16'h7869] = 8'hAD;
mem[16'h786A] = 8'hD0;
mem[16'h786B] = 8'h4D;
mem[16'h786C] = 8'h38;
mem[16'h786D] = 8'hED;
mem[16'h786E] = 8'h63;
mem[16'h786F] = 8'h79;
mem[16'h7870] = 8'h20;
mem[16'h7871] = 8'h62;
mem[16'h7872] = 8'h65;
mem[16'h7873] = 8'hC9;
mem[16'h7874] = 8'h04;
mem[16'h7875] = 8'hB0;
mem[16'h7876] = 8'h08;
mem[16'h7877] = 8'hA9;
mem[16'h7878] = 8'hC8;
mem[16'h7879] = 8'h20;
mem[16'h787A] = 8'hA8;
mem[16'h787B] = 8'hFC;
mem[16'h787C] = 8'h4C;
mem[16'h787D] = 8'h8E;
mem[16'h787E] = 8'h48;
mem[16'h787F] = 8'h20;
mem[16'h7880] = 8'h48;
mem[16'h7881] = 8'h79;
mem[16'h7882] = 8'hA9;
mem[16'h7883] = 8'h00;
mem[16'h7884] = 8'h8D;
mem[16'h7885] = 8'h33;
mem[16'h7886] = 8'h7B;
mem[16'h7887] = 8'hAD;
mem[16'h7888] = 8'hDF;
mem[16'h7889] = 8'h91;
mem[16'h788A] = 8'h8D;
mem[16'h788B] = 8'hDB;
mem[16'h788C] = 8'h91;
mem[16'h788D] = 8'h60;
mem[16'h788E] = 8'hAD;
mem[16'h788F] = 8'h62;
mem[16'h7890] = 8'h79;
mem[16'h7891] = 8'h38;
mem[16'h7892] = 8'hE9;
mem[16'h7893] = 8'h02;
mem[16'h7894] = 8'hC9;
mem[16'h7895] = 8'h05;
mem[16'h7896] = 8'h90;
mem[16'h7897] = 8'h15;
mem[16'h7898] = 8'h8D;
mem[16'h7899] = 8'h62;
mem[16'h789A] = 8'h79;
mem[16'h789B] = 8'h20;
mem[16'h789C] = 8'h16;
mem[16'h789D] = 8'h79;
mem[16'h789E] = 8'hAE;
mem[16'h789F] = 8'h34;
mem[16'h78A0] = 8'h7B;
mem[16'h78A1] = 8'hBD;
mem[16'h78A2] = 8'h2C;
mem[16'h78A3] = 8'h5F;
mem[16'h78A4] = 8'h18;
mem[16'h78A5] = 8'h69;
mem[16'h78A6] = 8'h0C;
mem[16'h78A7] = 8'h38;
mem[16'h78A8] = 8'hED;
mem[16'h78A9] = 8'h62;
mem[16'h78AA] = 8'h79;
mem[16'h78AB] = 8'h90;
mem[16'h78AC] = 8'h0F;
mem[16'h78AD] = 8'h20;
mem[16'h78AE] = 8'h7F;
mem[16'h78AF] = 8'h79;
mem[16'h78B0] = 8'hA9;
mem[16'h78B1] = 8'h00;
mem[16'h78B2] = 8'h8D;
mem[16'h78B3] = 8'h33;
mem[16'h78B4] = 8'h7B;
mem[16'h78B5] = 8'hAD;
mem[16'h78B6] = 8'hDF;
mem[16'h78B7] = 8'h91;
mem[16'h78B8] = 8'h8D;
mem[16'h78B9] = 8'hDB;
mem[16'h78BA] = 8'h91;
mem[16'h78BB] = 8'h60;
mem[16'h78BC] = 8'hAD;
mem[16'h78BD] = 8'hCF;
mem[16'h78BE] = 8'h4D;
mem[16'h78BF] = 8'h18;
mem[16'h78C0] = 8'h69;
mem[16'h78C1] = 8'h0E;
mem[16'h78C2] = 8'h38;
mem[16'h78C3] = 8'hED;
mem[16'h78C4] = 8'h62;
mem[16'h78C5] = 8'h79;
mem[16'h78C6] = 8'h20;
mem[16'h78C7] = 8'h62;
mem[16'h78C8] = 8'h65;
mem[16'h78C9] = 8'hC9;
mem[16'h78CA] = 8'h05;
mem[16'h78CB] = 8'hB0;
mem[16'h78CC] = 8'hEE;
mem[16'h78CD] = 8'hAD;
mem[16'h78CE] = 8'hD0;
mem[16'h78CF] = 8'h4D;
mem[16'h78D0] = 8'h38;
mem[16'h78D1] = 8'hED;
mem[16'h78D2] = 8'h63;
mem[16'h78D3] = 8'h79;
mem[16'h78D4] = 8'h20;
mem[16'h78D5] = 8'h62;
mem[16'h78D6] = 8'h65;
mem[16'h78D7] = 8'hC9;
mem[16'h78D8] = 8'h04;
mem[16'h78D9] = 8'hB0;
mem[16'h78DA] = 8'hE0;
mem[16'h78DB] = 8'hA9;
mem[16'h78DC] = 8'hC8;
mem[16'h78DD] = 8'h20;
mem[16'h78DE] = 8'hA8;
mem[16'h78DF] = 8'hFC;
mem[16'h78E0] = 8'h4C;
mem[16'h78E1] = 8'h8E;
mem[16'h78E2] = 8'h48;
mem[16'h78E3] = 8'hCE;
mem[16'h78E4] = 8'hAD;
mem[16'h78E5] = 8'h63;
mem[16'h78E6] = 8'h79;
mem[16'h78E7] = 8'h85;
mem[16'h78E8] = 8'h56;
mem[16'h78E9] = 8'hAC;
mem[16'h78EA] = 8'h62;
mem[16'h78EB] = 8'h79;
mem[16'h78EC] = 8'h84;
mem[16'h78ED] = 8'h57;
mem[16'h78EE] = 8'hB9;
mem[16'h78EF] = 8'h3E;
mem[16'h78F0] = 8'h8C;
mem[16'h78F1] = 8'hAA;
mem[16'h78F2] = 8'hBD;
mem[16'h78F3] = 8'h94;
mem[16'h78F4] = 8'h8E;
mem[16'h78F5] = 8'hAA;
mem[16'h78F6] = 8'hBD;
mem[16'h78F7] = 8'h08;
mem[16'h78F8] = 8'h79;
mem[16'h78F9] = 8'hBC;
mem[16'h78FA] = 8'h0F;
mem[16'h78FB] = 8'h79;
mem[16'h78FC] = 8'h20;
mem[16'h78FD] = 8'hD1;
mem[16'h78FE] = 8'h8A;
mem[16'h78FF] = 8'hA9;
mem[16'h7900] = 8'h24;
mem[16'h7901] = 8'h8D;
mem[16'h7902] = 8'hCA;
mem[16'h7903] = 8'h8A;
mem[16'h7904] = 8'h20;
mem[16'h7905] = 8'h79;
mem[16'h7906] = 8'h8A;
mem[16'h7907] = 8'h60;
mem[16'h7908] = 8'hBD;
mem[16'h7909] = 8'h99;
mem[16'h790A] = 8'h75;
mem[16'h790B] = 8'h51;
mem[16'h790C] = 8'h2D;
mem[16'h790D] = 8'h09;
mem[16'h790E] = 8'hE5;
mem[16'h790F] = 8'h95;
mem[16'h7910] = 8'h95;
mem[16'h7911] = 8'h95;
mem[16'h7912] = 8'h95;
mem[16'h7913] = 8'h95;
mem[16'h7914] = 8'h95;
mem[16'h7915] = 8'h94;
mem[16'h7916] = 8'hAD;
mem[16'h7917] = 8'h63;
mem[16'h7918] = 8'h79;
mem[16'h7919] = 8'h85;
mem[16'h791A] = 8'h56;
mem[16'h791B] = 8'hAC;
mem[16'h791C] = 8'h62;
mem[16'h791D] = 8'h79;
mem[16'h791E] = 8'h84;
mem[16'h791F] = 8'h57;
mem[16'h7920] = 8'hB9;
mem[16'h7921] = 8'h3E;
mem[16'h7922] = 8'h8C;
mem[16'h7923] = 8'hAA;
mem[16'h7924] = 8'hBD;
mem[16'h7925] = 8'h94;
mem[16'h7926] = 8'h8E;
mem[16'h7927] = 8'hAA;
mem[16'h7928] = 8'hBD;
mem[16'h7929] = 8'h3A;
mem[16'h792A] = 8'h79;
mem[16'h792B] = 8'hBC;
mem[16'h792C] = 8'h41;
mem[16'h792D] = 8'h79;
mem[16'h792E] = 8'h20;
mem[16'h792F] = 8'hD1;
mem[16'h7930] = 8'h8A;
mem[16'h7931] = 8'hA9;
mem[16'h7932] = 8'h24;
mem[16'h7933] = 8'h8D;
mem[16'h7934] = 8'hCA;
mem[16'h7935] = 8'h8A;
mem[16'h7936] = 8'h20;
mem[16'h7937] = 8'h79;
mem[16'h7938] = 8'h8A;
mem[16'h7939] = 8'h60;
mem[16'h793A] = 8'hC1;
mem[16'h793B] = 8'h9D;
mem[16'h793C] = 8'h79;
mem[16'h793D] = 8'h55;
mem[16'h793E] = 8'h31;
mem[16'h793F] = 8'h0D;
mem[16'h7940] = 8'hE9;
mem[16'h7941] = 8'h94;
mem[16'h7942] = 8'h94;
mem[16'h7943] = 8'h94;
mem[16'h7944] = 8'h94;
mem[16'h7945] = 8'h94;
mem[16'h7946] = 8'h94;
mem[16'h7947] = 8'h93;
mem[16'h7948] = 8'hA9;
mem[16'h7949] = 8'h64;
mem[16'h794A] = 8'hA0;
mem[16'h794B] = 8'h79;
mem[16'h794C] = 8'h20;
mem[16'h794D] = 8'h86;
mem[16'h794E] = 8'h68;
mem[16'h794F] = 8'hA9;
mem[16'h7950] = 8'h1B;
mem[16'h7951] = 8'h8D;
mem[16'h7952] = 8'h7F;
mem[16'h7953] = 8'h68;
mem[16'h7954] = 8'hAD;
mem[16'h7955] = 8'h62;
mem[16'h7956] = 8'h79;
mem[16'h7957] = 8'h85;
mem[16'h7958] = 8'h57;
mem[16'h7959] = 8'hAD;
mem[16'h795A] = 8'h63;
mem[16'h795B] = 8'h79;
mem[16'h795C] = 8'h85;
mem[16'h795D] = 8'h56;
mem[16'h795E] = 8'h20;
mem[16'h795F] = 8'hE6;
mem[16'h7960] = 8'h67;
mem[16'h7961] = 8'h60;
mem[16'h7962] = 8'h33;
mem[16'h7963] = 8'h30;
mem[16'h7964] = 8'h00;
mem[16'h7965] = 8'h28;
mem[16'h7966] = 8'h00;
mem[16'h7967] = 8'h00;
mem[16'h7968] = 8'h3A;
mem[16'h7969] = 8'h00;
mem[16'h796A] = 8'h00;
mem[16'h796B] = 8'h2A;
mem[16'h796C] = 8'h01;
mem[16'h796D] = 8'h40;
mem[16'h796E] = 8'h2A;
mem[16'h796F] = 8'h01;
mem[16'h7970] = 8'h40;
mem[16'h7971] = 8'h2A;
mem[16'h7972] = 8'h00;
mem[16'h7973] = 8'h40;
mem[16'h7974] = 8'h0A;
mem[16'h7975] = 8'h00;
mem[16'h7976] = 8'h50;
mem[16'h7977] = 8'h0A;
mem[16'h7978] = 8'h00;
mem[16'h7979] = 8'h54;
mem[16'h797A] = 8'h0A;
mem[16'h797B] = 8'h00;
mem[16'h797C] = 8'h55;
mem[16'h797D] = 8'h0A;
mem[16'h797E] = 8'h00;
mem[16'h797F] = 8'hA9;
mem[16'h7980] = 8'h99;
mem[16'h7981] = 8'hA0;
mem[16'h7982] = 8'h79;
mem[16'h7983] = 8'h20;
mem[16'h7984] = 8'h86;
mem[16'h7985] = 8'h68;
mem[16'h7986] = 8'hA9;
mem[16'h7987] = 8'h1B;
mem[16'h7988] = 8'h8D;
mem[16'h7989] = 8'h7F;
mem[16'h798A] = 8'h68;
mem[16'h798B] = 8'hAD;
mem[16'h798C] = 8'h62;
mem[16'h798D] = 8'h79;
mem[16'h798E] = 8'h85;
mem[16'h798F] = 8'h57;
mem[16'h7990] = 8'hAD;
mem[16'h7991] = 8'h63;
mem[16'h7992] = 8'h79;
mem[16'h7993] = 8'h85;
mem[16'h7994] = 8'h56;
mem[16'h7995] = 8'h20;
mem[16'h7996] = 8'hE6;
mem[16'h7997] = 8'h67;
mem[16'h7998] = 8'h60;
mem[16'h7999] = 8'h14;
mem[16'h799A] = 8'h00;
mem[16'h799B] = 8'h00;
mem[16'h799C] = 8'h5C;
mem[16'h799D] = 8'h00;
mem[16'h799E] = 8'h00;
mem[16'h799F] = 8'h55;
mem[16'h79A0] = 8'h00;
mem[16'h79A1] = 8'h00;
mem[16'h79A2] = 8'h55;
mem[16'h79A3] = 8'h02;
mem[16'h79A4] = 8'h00;
mem[16'h79A5] = 8'h54;
mem[16'h79A6] = 8'h02;
mem[16'h79A7] = 8'h00;
mem[16'h79A8] = 8'h50;
mem[16'h79A9] = 8'h02;
mem[16'h79AA] = 8'h00;
mem[16'h79AB] = 8'h50;
mem[16'h79AC] = 8'h0A;
mem[16'h79AD] = 8'h00;
mem[16'h79AE] = 8'h50;
mem[16'h79AF] = 8'h2A;
mem[16'h79B0] = 8'h00;
mem[16'h79B1] = 8'h50;
mem[16'h79B2] = 8'h2A;
mem[16'h79B3] = 8'h01;
mem[16'h79B4] = 8'hAD;
mem[16'h79B5] = 8'h33;
mem[16'h79B6] = 8'h7B;
mem[16'h79B7] = 8'hD0;
mem[16'h79B8] = 8'h5E;
mem[16'h79B9] = 8'hAD;
mem[16'h79BA] = 8'hCE;
mem[16'h79BB] = 8'h44;
mem[16'h79BC] = 8'hC9;
mem[16'h79BD] = 8'h04;
mem[16'h79BE] = 8'h90;
mem[16'h79BF] = 8'h03;
mem[16'h79C0] = 8'h4C;
mem[16'h79C1] = 8'h63;
mem[16'h79C2] = 8'h7A;
mem[16'h79C3] = 8'hA9;
mem[16'h79C4] = 8'h00;
mem[16'h79C5] = 8'h8D;
mem[16'h79C6] = 8'h35;
mem[16'h79C7] = 8'h7B;
mem[16'h79C8] = 8'hAD;
mem[16'h79C9] = 8'h13;
mem[16'h79CA] = 8'h87;
mem[16'h79CB] = 8'h29;
mem[16'h79CC] = 8'h03;
mem[16'h79CD] = 8'hC9;
mem[16'h79CE] = 8'h03;
mem[16'h79CF] = 8'h90;
mem[16'h79D0] = 8'h47;
mem[16'h79D1] = 8'hAD;
mem[16'h79D2] = 8'h35;
mem[16'h79D3] = 8'h7B;
mem[16'h79D4] = 8'hF0;
mem[16'h79D5] = 8'h01;
mem[16'h79D6] = 8'h60;
mem[16'h79D7] = 8'hA9;
mem[16'h79D8] = 8'h01;
mem[16'h79D9] = 8'h8D;
mem[16'h79DA] = 8'h35;
mem[16'h79DB] = 8'h7B;
mem[16'h79DC] = 8'hAD;
mem[16'h79DD] = 8'hB1;
mem[16'h79DE] = 8'h4A;
mem[16'h79DF] = 8'hF0;
mem[16'h79E0] = 8'h3B;
mem[16'h79E1] = 8'hAD;
mem[16'h79E2] = 8'h14;
mem[16'h79E3] = 8'h87;
mem[16'h79E4] = 8'h29;
mem[16'h79E5] = 8'h03;
mem[16'h79E6] = 8'hCD;
mem[16'h79E7] = 8'hB1;
mem[16'h79E8] = 8'h4A;
mem[16'h79E9] = 8'h90;
mem[16'h79EA] = 8'h02;
mem[16'h79EB] = 8'hA9;
mem[16'h79EC] = 8'h00;
mem[16'h79ED] = 8'hA8;
mem[16'h79EE] = 8'h8C;
mem[16'h79EF] = 8'h34;
mem[16'h79F0] = 8'h7B;
mem[16'h79F1] = 8'hAD;
mem[16'h79F2] = 8'h03;
mem[16'h79F3] = 8'h54;
mem[16'h79F4] = 8'h8D;
mem[16'h79F5] = 8'h63;
mem[16'h79F6] = 8'h79;
mem[16'h79F7] = 8'hB9;
mem[16'h79F8] = 8'h00;
mem[16'h79F9] = 8'h54;
mem[16'h79FA] = 8'hC9;
mem[16'h79FB] = 8'hF0;
mem[16'h79FC] = 8'hB0;
mem[16'h79FD] = 8'h1E;
mem[16'h79FE] = 8'h38;
mem[16'h79FF] = 8'hED;
mem[16'h7A00] = 8'h0C;
mem[16'h7A01] = 8'h54;
mem[16'h7A02] = 8'h90;
mem[16'h7A03] = 8'h13;
mem[16'h7A04] = 8'hE9;
mem[16'h7A05] = 8'h21;
mem[16'h7A06] = 8'h90;
mem[16'h7A07] = 8'h0F;
mem[16'h7A08] = 8'hC9;
mem[16'h7A09] = 8'hC8;
mem[16'h7A0A] = 8'hB0;
mem[16'h7A0B] = 8'h0B;
mem[16'h7A0C] = 8'h8D;
mem[16'h7A0D] = 8'h62;
mem[16'h7A0E] = 8'h79;
mem[16'h7A0F] = 8'h20;
mem[16'h7A10] = 8'h48;
mem[16'h7A11] = 8'h79;
mem[16'h7A12] = 8'hA9;
mem[16'h7A13] = 8'hFF;
mem[16'h7A14] = 8'h8D;
mem[16'h7A15] = 8'h33;
mem[16'h7A16] = 8'h7B;
mem[16'h7A17] = 8'h60;
mem[16'h7A18] = 8'hC9;
mem[16'h7A19] = 8'h01;
mem[16'h7A1A] = 8'h90;
mem[16'h7A1B] = 8'h20;
mem[16'h7A1C] = 8'hAD;
mem[16'h7A1D] = 8'h14;
mem[16'h7A1E] = 8'h87;
mem[16'h7A1F] = 8'h29;
mem[16'h7A20] = 8'h03;
mem[16'h7A21] = 8'hCD;
mem[16'h7A22] = 8'hB2;
mem[16'h7A23] = 8'h4A;
mem[16'h7A24] = 8'h90;
mem[16'h7A25] = 8'h02;
mem[16'h7A26] = 8'hA9;
mem[16'h7A27] = 8'h00;
mem[16'h7A28] = 8'hA8;
mem[16'h7A29] = 8'h8C;
mem[16'h7A2A] = 8'h34;
mem[16'h7A2B] = 8'h7B;
mem[16'h7A2C] = 8'hAD;
mem[16'h7A2D] = 8'h13;
mem[16'h7A2E] = 8'h51;
mem[16'h7A2F] = 8'h8D;
mem[16'h7A30] = 8'h63;
mem[16'h7A31] = 8'h79;
mem[16'h7A32] = 8'hB9;
mem[16'h7A33] = 8'h10;
mem[16'h7A34] = 8'h51;
mem[16'h7A35] = 8'h38;
mem[16'h7A36] = 8'hED;
mem[16'h7A37] = 8'h1F;
mem[16'h7A38] = 8'h51;
mem[16'h7A39] = 8'h4C;
mem[16'h7A3A] = 8'h02;
mem[16'h7A3B] = 8'h7A;
mem[16'h7A3C] = 8'hAD;
mem[16'h7A3D] = 8'h14;
mem[16'h7A3E] = 8'h87;
mem[16'h7A3F] = 8'h29;
mem[16'h7A40] = 8'h03;
mem[16'h7A41] = 8'hCD;
mem[16'h7A42] = 8'hB3;
mem[16'h7A43] = 8'h4A;
mem[16'h7A44] = 8'h90;
mem[16'h7A45] = 8'h02;
mem[16'h7A46] = 8'hA9;
mem[16'h7A47] = 8'h00;
mem[16'h7A48] = 8'hA8;
mem[16'h7A49] = 8'h8C;
mem[16'h7A4A] = 8'h34;
mem[16'h7A4B] = 8'h7B;
mem[16'h7A4C] = 8'hAD;
mem[16'h7A4D] = 8'h23;
mem[16'h7A4E] = 8'h53;
mem[16'h7A4F] = 8'h8D;
mem[16'h7A50] = 8'h63;
mem[16'h7A51] = 8'h79;
mem[16'h7A52] = 8'hB9;
mem[16'h7A53] = 8'h1F;
mem[16'h7A54] = 8'h53;
mem[16'h7A55] = 8'hC9;
mem[16'h7A56] = 8'hF0;
mem[16'h7A57] = 8'h90;
mem[16'h7A58] = 8'h03;
mem[16'h7A59] = 8'h4C;
mem[16'h7A5A] = 8'hD1;
mem[16'h7A5B] = 8'h79;
mem[16'h7A5C] = 8'h38;
mem[16'h7A5D] = 8'hED;
mem[16'h7A5E] = 8'h27;
mem[16'h7A5F] = 8'h53;
mem[16'h7A60] = 8'h4C;
mem[16'h7A61] = 8'h02;
mem[16'h7A62] = 8'h7A;
mem[16'h7A63] = 8'hAD;
mem[16'h7A64] = 8'h13;
mem[16'h7A65] = 8'h87;
mem[16'h7A66] = 8'h29;
mem[16'h7A67] = 8'h07;
mem[16'h7A68] = 8'hC9;
mem[16'h7A69] = 8'h07;
mem[16'h7A6A] = 8'h90;
mem[16'h7A6B] = 8'h3C;
mem[16'h7A6C] = 8'hAD;
mem[16'h7A6D] = 8'hB1;
mem[16'h7A6E] = 8'h4A;
mem[16'h7A6F] = 8'hF0;
mem[16'h7A70] = 8'h36;
mem[16'h7A71] = 8'hAD;
mem[16'h7A72] = 8'h14;
mem[16'h7A73] = 8'h87;
mem[16'h7A74] = 8'h29;
mem[16'h7A75] = 8'h03;
mem[16'h7A76] = 8'hCD;
mem[16'h7A77] = 8'hB1;
mem[16'h7A78] = 8'h4A;
mem[16'h7A79] = 8'h90;
mem[16'h7A7A] = 8'h02;
mem[16'h7A7B] = 8'hA9;
mem[16'h7A7C] = 8'h00;
mem[16'h7A7D] = 8'hA8;
mem[16'h7A7E] = 8'h8C;
mem[16'h7A7F] = 8'h34;
mem[16'h7A80] = 8'h7B;
mem[16'h7A81] = 8'hAD;
mem[16'h7A82] = 8'h03;
mem[16'h7A83] = 8'h54;
mem[16'h7A84] = 8'h8D;
mem[16'h7A85] = 8'h63;
mem[16'h7A86] = 8'h79;
mem[16'h7A87] = 8'hB9;
mem[16'h7A88] = 8'h00;
mem[16'h7A89] = 8'h54;
mem[16'h7A8A] = 8'hC9;
mem[16'h7A8B] = 8'hF0;
mem[16'h7A8C] = 8'hB0;
mem[16'h7A8D] = 8'h19;
mem[16'h7A8E] = 8'h38;
mem[16'h7A8F] = 8'hED;
mem[16'h7A90] = 8'h0C;
mem[16'h7A91] = 8'h54;
mem[16'h7A92] = 8'h90;
mem[16'h7A93] = 8'h13;
mem[16'h7A94] = 8'hE9;
mem[16'h7A95] = 8'h21;
mem[16'h7A96] = 8'h90;
mem[16'h7A97] = 8'h0F;
mem[16'h7A98] = 8'hC9;
mem[16'h7A99] = 8'hC8;
mem[16'h7A9A] = 8'hB0;
mem[16'h7A9B] = 8'h0B;
mem[16'h7A9C] = 8'h8D;
mem[16'h7A9D] = 8'h62;
mem[16'h7A9E] = 8'h79;
mem[16'h7A9F] = 8'h20;
mem[16'h7AA0] = 8'h48;
mem[16'h7AA1] = 8'h79;
mem[16'h7AA2] = 8'hA9;
mem[16'h7AA3] = 8'hFF;
mem[16'h7AA4] = 8'h8D;
mem[16'h7AA5] = 8'h33;
mem[16'h7AA6] = 8'h7B;
mem[16'h7AA7] = 8'h60;
mem[16'h7AA8] = 8'hC9;
mem[16'h7AA9] = 8'h05;
mem[16'h7AAA] = 8'h90;
mem[16'h7AAB] = 8'h20;
mem[16'h7AAC] = 8'hAD;
mem[16'h7AAD] = 8'h14;
mem[16'h7AAE] = 8'h87;
mem[16'h7AAF] = 8'h29;
mem[16'h7AB0] = 8'h03;
mem[16'h7AB1] = 8'hCD;
mem[16'h7AB2] = 8'hB2;
mem[16'h7AB3] = 8'h4A;
mem[16'h7AB4] = 8'h90;
mem[16'h7AB5] = 8'h02;
mem[16'h7AB6] = 8'hA9;
mem[16'h7AB7] = 8'h00;
mem[16'h7AB8] = 8'hA8;
mem[16'h7AB9] = 8'h8C;
mem[16'h7ABA] = 8'h34;
mem[16'h7ABB] = 8'h7B;
mem[16'h7ABC] = 8'hAD;
mem[16'h7ABD] = 8'h13;
mem[16'h7ABE] = 8'h51;
mem[16'h7ABF] = 8'h8D;
mem[16'h7AC0] = 8'h63;
mem[16'h7AC1] = 8'h79;
mem[16'h7AC2] = 8'hB9;
mem[16'h7AC3] = 8'h10;
mem[16'h7AC4] = 8'h51;
mem[16'h7AC5] = 8'h38;
mem[16'h7AC6] = 8'hED;
mem[16'h7AC7] = 8'h1F;
mem[16'h7AC8] = 8'h51;
mem[16'h7AC9] = 8'h4C;
mem[16'h7ACA] = 8'h92;
mem[16'h7ACB] = 8'h7A;
mem[16'h7ACC] = 8'hC9;
mem[16'h7ACD] = 8'h04;
mem[16'h7ACE] = 8'h90;
mem[16'h7ACF] = 8'h24;
mem[16'h7AD0] = 8'hAD;
mem[16'h7AD1] = 8'h14;
mem[16'h7AD2] = 8'h87;
mem[16'h7AD3] = 8'h29;
mem[16'h7AD4] = 8'h03;
mem[16'h7AD5] = 8'hCD;
mem[16'h7AD6] = 8'hB3;
mem[16'h7AD7] = 8'h4A;
mem[16'h7AD8] = 8'h90;
mem[16'h7AD9] = 8'h02;
mem[16'h7ADA] = 8'hA9;
mem[16'h7ADB] = 8'h00;
mem[16'h7ADC] = 8'hA8;
mem[16'h7ADD] = 8'h8C;
mem[16'h7ADE] = 8'h34;
mem[16'h7ADF] = 8'h7B;
mem[16'h7AE0] = 8'hAD;
mem[16'h7AE1] = 8'h23;
mem[16'h7AE2] = 8'h53;
mem[16'h7AE3] = 8'h8D;
mem[16'h7AE4] = 8'h63;
mem[16'h7AE5] = 8'h79;
mem[16'h7AE6] = 8'hB9;
mem[16'h7AE7] = 8'h1F;
mem[16'h7AE8] = 8'h53;
mem[16'h7AE9] = 8'hC9;
mem[16'h7AEA] = 8'hF0;
mem[16'h7AEB] = 8'hB0;
mem[16'h7AEC] = 8'hBA;
mem[16'h7AED] = 8'h38;
mem[16'h7AEE] = 8'hED;
mem[16'h7AEF] = 8'h27;
mem[16'h7AF0] = 8'h53;
mem[16'h7AF1] = 8'h4C;
mem[16'h7AF2] = 8'h92;
mem[16'h7AF3] = 8'h7A;
mem[16'h7AF4] = 8'hC9;
mem[16'h7AF5] = 8'h02;
mem[16'h7AF6] = 8'h90;
mem[16'h7AF7] = 8'h32;
mem[16'h7AF8] = 8'hAD;
mem[16'h7AF9] = 8'h14;
mem[16'h7AFA] = 8'h87;
mem[16'h7AFB] = 8'h29;
mem[16'h7AFC] = 8'h04;
mem[16'h7AFD] = 8'hCD;
mem[16'h7AFE] = 8'hAF;
mem[16'h7AFF] = 8'h4A;
mem[16'h7B00] = 8'h90;
mem[16'h7B01] = 8'h02;
mem[16'h7B02] = 8'hA9;
mem[16'h7B03] = 8'h00;
mem[16'h7B04] = 8'hA8;
mem[16'h7B05] = 8'h8C;
mem[16'h7B06] = 8'h34;
mem[16'h7B07] = 8'h7B;
mem[16'h7B08] = 8'hB9;
mem[16'h7B09] = 8'h1E;
mem[16'h7B0A] = 8'h5F;
mem[16'h7B0B] = 8'h8D;
mem[16'h7B0C] = 8'h63;
mem[16'h7B0D] = 8'h79;
mem[16'h7B0E] = 8'hB9;
mem[16'h7B0F] = 8'h2C;
mem[16'h7B10] = 8'h5F;
mem[16'h7B11] = 8'hC9;
mem[16'h7B12] = 8'h14;
mem[16'h7B13] = 8'h90;
mem[16'h7B14] = 8'h14;
mem[16'h7B15] = 8'h18;
mem[16'h7B16] = 8'h69;
mem[16'h7B17] = 8'h1F;
mem[16'h7B18] = 8'hB0;
mem[16'h7B19] = 8'h0F;
mem[16'h7B1A] = 8'hC9;
mem[16'h7B1B] = 8'hDC;
mem[16'h7B1C] = 8'hB0;
mem[16'h7B1D] = 8'h0B;
mem[16'h7B1E] = 8'h8D;
mem[16'h7B1F] = 8'h62;
mem[16'h7B20] = 8'h79;
mem[16'h7B21] = 8'h20;
mem[16'h7B22] = 8'h7F;
mem[16'h7B23] = 8'h79;
mem[16'h7B24] = 8'hA9;
mem[16'h7B25] = 8'hFF;
mem[16'h7B26] = 8'h8D;
mem[16'h7B27] = 8'h33;
mem[16'h7B28] = 8'h7B;
mem[16'h7B29] = 8'h60;
mem[16'h7B2A] = 8'hA9;
mem[16'h7B2B] = 8'h08;
mem[16'h7B2C] = 8'hA8;
mem[16'h7B2D] = 8'h8C;
mem[16'h7B2E] = 8'h34;
mem[16'h7B2F] = 8'h7B;
mem[16'h7B30] = 8'h4C;
mem[16'h7B31] = 8'h08;
mem[16'h7B32] = 8'h7B;
mem[16'h7B33] = 8'h00;
mem[16'h7B34] = 8'h54;
mem[16'h7B35] = 8'h00;
mem[16'h7B36] = 8'hAD;
mem[16'h7B37] = 8'h5A;
mem[16'h7B38] = 8'h74;
mem[16'h7B39] = 8'hD0;
mem[16'h7B3A] = 8'h01;
mem[16'h7B3B] = 8'h60;
mem[16'h7B3C] = 8'hA9;
mem[16'h7B3D] = 8'hCD;
mem[16'h7B3E] = 8'h8D;
mem[16'h7B3F] = 8'h84;
mem[16'h7B40] = 8'h7B;
mem[16'h7B41] = 8'hA9;
mem[16'h7B42] = 8'h17;
mem[16'h7B43] = 8'h8D;
mem[16'h7B44] = 8'h87;
mem[16'h7B45] = 8'h7B;
mem[16'h7B46] = 8'h8D;
mem[16'h7B47] = 8'h88;
mem[16'h7B48] = 8'h7B;
mem[16'h7B49] = 8'h8D;
mem[16'h7B4A] = 8'h89;
mem[16'h7B4B] = 8'h7B;
mem[16'h7B4C] = 8'hA9;
mem[16'h7B4D] = 8'h1E;
mem[16'h7B4E] = 8'h8D;
mem[16'h7B4F] = 8'h92;
mem[16'h7B50] = 8'h73;
mem[16'h7B51] = 8'hA2;
mem[16'h7B52] = 8'h00;
mem[16'h7B53] = 8'h86;
mem[16'h7B54] = 8'h70;
mem[16'h7B55] = 8'h20;
mem[16'h7B56] = 8'h8A;
mem[16'h7B57] = 8'h7B;
mem[16'h7B58] = 8'hAD;
mem[16'h7B59] = 8'h5A;
mem[16'h7B5A] = 8'h74;
mem[16'h7B5B] = 8'hC9;
mem[16'h7B5C] = 8'h02;
mem[16'h7B5D] = 8'h90;
mem[16'h7B5E] = 8'h1F;
mem[16'h7B5F] = 8'hA9;
mem[16'h7B60] = 8'h7D;
mem[16'h7B61] = 8'h8D;
mem[16'h7B62] = 8'h85;
mem[16'h7B63] = 8'h7B;
mem[16'h7B64] = 8'hA2;
mem[16'h7B65] = 8'h01;
mem[16'h7B66] = 8'h86;
mem[16'h7B67] = 8'h70;
mem[16'h7B68] = 8'h20;
mem[16'h7B69] = 8'h8A;
mem[16'h7B6A] = 8'h7B;
mem[16'h7B6B] = 8'hAD;
mem[16'h7B6C] = 8'h5A;
mem[16'h7B6D] = 8'h74;
mem[16'h7B6E] = 8'hC9;
mem[16'h7B6F] = 8'h03;
mem[16'h7B70] = 8'h90;
mem[16'h7B71] = 8'h0C;
mem[16'h7B72] = 8'hA9;
mem[16'h7B73] = 8'h2D;
mem[16'h7B74] = 8'h8D;
mem[16'h7B75] = 8'h86;
mem[16'h7B76] = 8'h7B;
mem[16'h7B77] = 8'hA2;
mem[16'h7B78] = 8'h02;
mem[16'h7B79] = 8'h86;
mem[16'h7B7A] = 8'h70;
mem[16'h7B7B] = 8'h20;
mem[16'h7B7C] = 8'h8A;
mem[16'h7B7D] = 8'h7B;
mem[16'h7B7E] = 8'hA9;
mem[16'h7B7F] = 8'h00;
mem[16'h7B80] = 8'h8D;
mem[16'h7B81] = 8'h93;
mem[16'h7B82] = 8'h73;
mem[16'h7B83] = 8'h60;
mem[16'h7B84] = 8'h41;
mem[16'h7B85] = 8'h4C;
mem[16'h7B86] = 8'h4C;
mem[16'h7B87] = 8'h31;
mem[16'h7B88] = 8'h0D;
mem[16'h7B89] = 8'h03;
mem[16'h7B8A] = 8'hA9;
mem[16'h7B8B] = 8'h10;
mem[16'h7B8C] = 8'hA0;
mem[16'h7B8D] = 8'h7C;
mem[16'h7B8E] = 8'h20;
mem[16'h7B8F] = 8'h86;
mem[16'h7B90] = 8'h68;
mem[16'h7B91] = 8'hA9;
mem[16'h7B92] = 8'h12;
mem[16'h7B93] = 8'h8D;
mem[16'h7B94] = 8'h7F;
mem[16'h7B95] = 8'h68;
mem[16'h7B96] = 8'hA6;
mem[16'h7B97] = 8'h70;
mem[16'h7B98] = 8'hBD;
mem[16'h7B99] = 8'h84;
mem[16'h7B9A] = 8'h7B;
mem[16'h7B9B] = 8'h85;
mem[16'h7B9C] = 8'h57;
mem[16'h7B9D] = 8'hBD;
mem[16'h7B9E] = 8'h87;
mem[16'h7B9F] = 8'h7B;
mem[16'h7BA0] = 8'h18;
mem[16'h7BA1] = 8'h69;
mem[16'h7BA2] = 8'h04;
mem[16'h7BA3] = 8'h85;
mem[16'h7BA4] = 8'h56;
mem[16'h7BA5] = 8'h20;
mem[16'h7BA6] = 8'hE6;
mem[16'h7BA7] = 8'h67;
mem[16'h7BA8] = 8'hA9;
mem[16'h7BA9] = 8'h22;
mem[16'h7BAA] = 8'hA0;
mem[16'h7BAB] = 8'h7C;
mem[16'h7BAC] = 8'h20;
mem[16'h7BAD] = 8'h2B;
mem[16'h7BAE] = 8'h8C;
mem[16'h7BAF] = 8'hA9;
mem[16'h7BB0] = 8'h10;
mem[16'h7BB1] = 8'h8D;
mem[16'h7BB2] = 8'h24;
mem[16'h7BB3] = 8'h8C;
mem[16'h7BB4] = 8'hA6;
mem[16'h7BB5] = 8'h70;
mem[16'h7BB6] = 8'hBD;
mem[16'h7BB7] = 8'h84;
mem[16'h7BB8] = 8'h7B;
mem[16'h7BB9] = 8'h18;
mem[16'h7BBA] = 8'h69;
mem[16'h7BBB] = 8'h15;
mem[16'h7BBC] = 8'h85;
mem[16'h7BBD] = 8'h57;
mem[16'h7BBE] = 8'hBD;
mem[16'h7BBF] = 8'h87;
mem[16'h7BC0] = 8'h7B;
mem[16'h7BC1] = 8'h18;
mem[16'h7BC2] = 8'h69;
mem[16'h7BC3] = 8'h02;
mem[16'h7BC4] = 8'h85;
mem[16'h7BC5] = 8'h56;
mem[16'h7BC6] = 8'h20;
mem[16'h7BC7] = 8'hA8;
mem[16'h7BC8] = 8'h8B;
mem[16'h7BC9] = 8'hAD;
mem[16'h7BCA] = 8'h0F;
mem[16'h7BCB] = 8'h7C;
mem[16'h7BCC] = 8'hF0;
mem[16'h7BCD] = 8'h1F;
mem[16'h7BCE] = 8'hA9;
mem[16'h7BCF] = 8'h32;
mem[16'h7BD0] = 8'hA0;
mem[16'h7BD1] = 8'h7C;
mem[16'h7BD2] = 8'h20;
mem[16'h7BD3] = 8'h2B;
mem[16'h7BD4] = 8'h8C;
mem[16'h7BD5] = 8'hA6;
mem[16'h7BD6] = 8'h70;
mem[16'h7BD7] = 8'hBD;
mem[16'h7BD8] = 8'h84;
mem[16'h7BD9] = 8'h7B;
mem[16'h7BDA] = 8'h18;
mem[16'h7BDB] = 8'h69;
mem[16'h7BDC] = 8'h23;
mem[16'h7BDD] = 8'h85;
mem[16'h7BDE] = 8'h57;
mem[16'h7BDF] = 8'hBD;
mem[16'h7BE0] = 8'h87;
mem[16'h7BE1] = 8'h7B;
mem[16'h7BE2] = 8'h85;
mem[16'h7BE3] = 8'h56;
mem[16'h7BE4] = 8'hA9;
mem[16'h7BE5] = 8'h14;
mem[16'h7BE6] = 8'h8D;
mem[16'h7BE7] = 8'h24;
mem[16'h7BE8] = 8'h8C;
mem[16'h7BE9] = 8'h20;
mem[16'h7BEA] = 8'hA8;
mem[16'h7BEB] = 8'h8B;
mem[16'h7BEC] = 8'h60;
mem[16'h7BED] = 8'hA9;
mem[16'h7BEE] = 8'h46;
mem[16'h7BEF] = 8'hA0;
mem[16'h7BF0] = 8'h7C;
mem[16'h7BF1] = 8'h20;
mem[16'h7BF2] = 8'h2B;
mem[16'h7BF3] = 8'h8C;
mem[16'h7BF4] = 8'hA6;
mem[16'h7BF5] = 8'h70;
mem[16'h7BF6] = 8'hBD;
mem[16'h7BF7] = 8'h84;
mem[16'h7BF8] = 8'h7B;
mem[16'h7BF9] = 8'h18;
mem[16'h7BFA] = 8'h69;
mem[16'h7BFB] = 8'h23;
mem[16'h7BFC] = 8'h85;
mem[16'h7BFD] = 8'h57;
mem[16'h7BFE] = 8'hBD;
mem[16'h7BFF] = 8'h87;
mem[16'h7C00] = 8'h7B;
mem[16'h7C01] = 8'h18;
mem[16'h7C02] = 8'h69;
mem[16'h7C03] = 8'h02;
mem[16'h7C04] = 8'h85;
mem[16'h7C05] = 8'h56;
mem[16'h7C06] = 8'hA9;
mem[16'h7C07] = 8'h10;
mem[16'h7C08] = 8'h8D;
mem[16'h7C09] = 8'h24;
mem[16'h7C0A] = 8'h8C;
mem[16'h7C0B] = 8'h20;
mem[16'h7C0C] = 8'hA8;
mem[16'h7C0D] = 8'h8B;
mem[16'h7C0E] = 8'h60;
mem[16'h7C0F] = 8'h01;
mem[16'h7C10] = 8'h00;
mem[16'h7C11] = 8'h00;
mem[16'h7C12] = 8'h40;
mem[16'h7C13] = 8'h00;
mem[16'h7C14] = 8'h00;
mem[16'h7C15] = 8'h7F;
mem[16'h7C16] = 8'h00;
mem[16'h7C17] = 8'h7E;
mem[16'h7C18] = 8'h7F;
mem[16'h7C19] = 8'h7F;
mem[16'h7C1A] = 8'h7F;
mem[16'h7C1B] = 8'h7F;
mem[16'h7C1C] = 8'h7C;
mem[16'h7C1D] = 8'h7F;
mem[16'h7C1E] = 8'h7F;
mem[16'h7C1F] = 8'h00;
mem[16'h7C20] = 8'h78;
mem[16'h7C21] = 8'h7F;
mem[16'h7C22] = 8'h00;
mem[16'h7C23] = 8'h70;
mem[16'h7C24] = 8'h00;
mem[16'h7C25] = 8'h7F;
mem[16'h7C26] = 8'h7F;
mem[16'h7C27] = 8'h7F;
mem[16'h7C28] = 8'h7F;
mem[16'h7C29] = 8'h7F;
mem[16'h7C2A] = 8'h7F;
mem[16'h7C2B] = 8'h7F;
mem[16'h7C2C] = 8'h7F;
mem[16'h7C2D] = 8'h7F;
mem[16'h7C2E] = 8'h7F;
mem[16'h7C2F] = 8'h7F;
mem[16'h7C30] = 8'h7F;
mem[16'h7C31] = 8'h7F;
mem[16'h7C32] = 8'h00;
mem[16'h7C33] = 8'h10;
mem[16'h7C34] = 8'h00;
mem[16'h7C35] = 8'h1C;
mem[16'h7C36] = 8'h03;
mem[16'h7C37] = 8'h17;
mem[16'h7C38] = 8'h7F;
mem[16'h7C39] = 8'h17;
mem[16'h7C3A] = 8'h7D;
mem[16'h7C3B] = 8'h05;
mem[16'h7C3C] = 8'h3F;
mem[16'h7C3D] = 8'h04;
mem[16'h7C3E] = 8'h0F;
mem[16'h7C3F] = 8'h11;
mem[16'h7C40] = 8'h0B;
mem[16'h7C41] = 8'h11;
mem[16'h7C42] = 8'h7F;
mem[16'h7C43] = 8'h1F;
mem[16'h7C44] = 8'h7F;
mem[16'h7C45] = 8'h07;
mem[16'h7C46] = 8'h03;
mem[16'h7C47] = 8'h00;
mem[16'h7C48] = 8'h0F;
mem[16'h7C49] = 8'h00;
mem[16'h7C4A] = 8'h0D;
mem[16'h7C4B] = 8'h00;
mem[16'h7C4C] = 8'h3F;
mem[16'h7C4D] = 8'h00;
mem[16'h7C4E] = 8'h7F;
mem[16'h7C4F] = 8'h7F;
mem[16'h7C50] = 8'h2F;
mem[16'h7C51] = 8'h55;
mem[16'h7C52] = 8'h7F;
mem[16'h7C53] = 8'h7F;
mem[16'h7C54] = 8'h7F;
mem[16'h7C55] = 8'h1F;
mem[16'h7C56] = 8'h00;
mem[16'h7C57] = 8'h50;
mem[16'h7C58] = 8'h02;
mem[16'h7C59] = 8'h00;
mem[16'h7C5A] = 8'h00;
mem[16'h7C5B] = 8'h50;
mem[16'h7C5C] = 8'h28;
mem[16'h7C5D] = 8'h01;
mem[16'h7C5E] = 8'h00;
mem[16'h7C5F] = 8'h30;
mem[16'h7C60] = 8'h24;
mem[16'h7C61] = 8'h00;
mem[16'h7C62] = 8'h00;
mem[16'h7C63] = 8'h06;
mem[16'h7C64] = 8'h30;
mem[16'h7C65] = 8'h00;
mem[16'h7C66] = 8'h40;
mem[16'h7C67] = 8'h38;
mem[16'h7C68] = 8'h40;
mem[16'h7C69] = 8'h01;
mem[16'h7C6A] = 8'h40;
mem[16'h7C6B] = 8'h38;
mem[16'h7C6C] = 8'h40;
mem[16'h7C6D] = 8'h01;
mem[16'h7C6E] = 8'h40;
mem[16'h7C6F] = 8'h38;
mem[16'h7C70] = 8'h40;
mem[16'h7C71] = 8'h01;
mem[16'h7C72] = 8'h00;
mem[16'h7C73] = 8'h06;
mem[16'h7C74] = 8'h30;
mem[16'h7C75] = 8'h00;
mem[16'h7C76] = 8'h00;
mem[16'h7C77] = 8'h30;
mem[16'h7C78] = 8'h24;
mem[16'h7C79] = 8'h00;
mem[16'h7C7A] = 8'h00;
mem[16'h7C7B] = 8'h50;
mem[16'h7C7C] = 8'h28;
mem[16'h7C7D] = 8'h01;
mem[16'h7C7E] = 8'h00;
mem[16'h7C7F] = 8'h50;
mem[16'h7C80] = 8'h02;
mem[16'h7C81] = 8'h00;
mem[16'h7C82] = 8'h00;
mem[16'h7C83] = 8'h28;
mem[16'h7C84] = 8'h01;
mem[16'h7C85] = 8'h00;
mem[16'h7C86] = 8'h00;
mem[16'h7C87] = 8'h28;
mem[16'h7C88] = 8'h54;
mem[16'h7C89] = 8'h00;
mem[16'h7C8A] = 8'h00;
mem[16'h7C8B] = 8'h18;
mem[16'h7C8C] = 8'h12;
mem[16'h7C8D] = 8'h00;
mem[16'h7C8E] = 8'h00;
mem[16'h7C8F] = 8'h03;
mem[16'h7C90] = 8'h18;
mem[16'h7C91] = 8'h00;
mem[16'h7C92] = 8'h20;
mem[16'h7C93] = 8'h1C;
mem[16'h7C94] = 8'h60;
mem[16'h7C95] = 8'h00;
mem[16'h7C96] = 8'h20;
mem[16'h7C97] = 8'h1C;
mem[16'h7C98] = 8'h60;
mem[16'h7C99] = 8'h00;
mem[16'h7C9A] = 8'h20;
mem[16'h7C9B] = 8'h1C;
mem[16'h7C9C] = 8'h60;
mem[16'h7C9D] = 8'h00;
mem[16'h7C9E] = 8'h00;
mem[16'h7C9F] = 8'h03;
mem[16'h7CA0] = 8'h18;
mem[16'h7CA1] = 8'h00;
mem[16'h7CA2] = 8'h00;
mem[16'h7CA3] = 8'h18;
mem[16'h7CA4] = 8'h12;
mem[16'h7CA5] = 8'h00;
mem[16'h7CA6] = 8'h00;
mem[16'h7CA7] = 8'h28;
mem[16'h7CA8] = 8'h54;
mem[16'h7CA9] = 8'h00;
mem[16'h7CAA] = 8'h00;
mem[16'h7CAB] = 8'h28;
mem[16'h7CAC] = 8'h01;
mem[16'h7CAD] = 8'h00;
mem[16'h7CAE] = 8'h00;
mem[16'h7CAF] = 8'h54;
mem[16'h7CB0] = 8'h00;
mem[16'h7CB1] = 8'h00;
mem[16'h7CB2] = 8'h00;
mem[16'h7CB3] = 8'h14;
mem[16'h7CB4] = 8'h2A;
mem[16'h7CB5] = 8'h00;
mem[16'h7CB6] = 8'h00;
mem[16'h7CB7] = 8'h0C;
mem[16'h7CB8] = 8'h09;
mem[16'h7CB9] = 8'h00;
mem[16'h7CBA] = 8'h40;
mem[16'h7CBB] = 8'h01;
mem[16'h7CBC] = 8'h0C;
mem[16'h7CBD] = 8'h00;
mem[16'h7CBE] = 8'h10;
mem[16'h7CBF] = 8'h0E;
mem[16'h7CC0] = 8'h30;
mem[16'h7CC1] = 8'h00;
mem[16'h7CC2] = 8'h10;
mem[16'h7CC3] = 8'h0E;
mem[16'h7CC4] = 8'h30;
mem[16'h7CC5] = 8'h00;
mem[16'h7CC6] = 8'h10;
mem[16'h7CC7] = 8'h0E;
mem[16'h7CC8] = 8'h30;
mem[16'h7CC9] = 8'h00;
mem[16'h7CCA] = 8'h40;
mem[16'h7CCB] = 8'h01;
mem[16'h7CCC] = 8'h0C;
mem[16'h7CCD] = 8'h00;
mem[16'h7CCE] = 8'h00;
mem[16'h7CCF] = 8'h0C;
mem[16'h7CD0] = 8'h09;
mem[16'h7CD1] = 8'h00;
mem[16'h7CD2] = 8'h00;
mem[16'h7CD3] = 8'h14;
mem[16'h7CD4] = 8'h2A;
mem[16'h7CD5] = 8'h00;
mem[16'h7CD6] = 8'h00;
mem[16'h7CD7] = 8'h54;
mem[16'h7CD8] = 8'h00;
mem[16'h7CD9] = 8'h00;
mem[16'h7CDA] = 8'h00;
mem[16'h7CDB] = 8'h2A;
mem[16'h7CDC] = 8'h00;
mem[16'h7CDD] = 8'h00;
mem[16'h7CDE] = 8'h00;
mem[16'h7CDF] = 8'h0A;
mem[16'h7CE0] = 8'h15;
mem[16'h7CE1] = 8'h00;
mem[16'h7CE2] = 8'h00;
mem[16'h7CE3] = 8'h46;
mem[16'h7CE4] = 8'h04;
mem[16'h7CE5] = 8'h00;
mem[16'h7CE6] = 8'h60;
mem[16'h7CE7] = 8'h00;
mem[16'h7CE8] = 8'h06;
mem[16'h7CE9] = 8'h00;
mem[16'h7CEA] = 8'h08;
mem[16'h7CEB] = 8'h07;
mem[16'h7CEC] = 8'h18;
mem[16'h7CED] = 8'h00;
mem[16'h7CEE] = 8'h08;
mem[16'h7CEF] = 8'h07;
mem[16'h7CF0] = 8'h18;
mem[16'h7CF1] = 8'h00;
mem[16'h7CF2] = 8'h08;
mem[16'h7CF3] = 8'h07;
mem[16'h7CF4] = 8'h18;
mem[16'h7CF5] = 8'h00;
mem[16'h7CF6] = 8'h60;
mem[16'h7CF7] = 8'h00;
mem[16'h7CF8] = 8'h06;
mem[16'h7CF9] = 8'h00;
mem[16'h7CFA] = 8'h00;
mem[16'h7CFB] = 8'h46;
mem[16'h7CFC] = 8'h04;
mem[16'h7CFD] = 8'h00;
mem[16'h7CFE] = 8'h00;
mem[16'h7CFF] = 8'h0A;
mem[16'h7D00] = 8'h15;
mem[16'h7D01] = 8'h00;
mem[16'h7D02] = 8'h00;
mem[16'h7D03] = 8'h2A;
mem[16'h7D04] = 8'h00;
mem[16'h7D05] = 8'h00;
mem[16'h7D06] = 8'h00;
mem[16'h7D07] = 8'h15;
mem[16'h7D08] = 8'h00;
mem[16'h7D09] = 8'h00;
mem[16'h7D0A] = 8'h00;
mem[16'h7D0B] = 8'h45;
mem[16'h7D0C] = 8'h0A;
mem[16'h7D0D] = 8'h00;
mem[16'h7D0E] = 8'h00;
mem[16'h7D0F] = 8'h23;
mem[16'h7D10] = 8'h02;
mem[16'h7D11] = 8'h00;
mem[16'h7D12] = 8'h30;
mem[16'h7D13] = 8'h00;
mem[16'h7D14] = 8'h03;
mem[16'h7D15] = 8'h00;
mem[16'h7D16] = 8'h44;
mem[16'h7D17] = 8'h03;
mem[16'h7D18] = 8'h0C;
mem[16'h7D19] = 8'h00;
mem[16'h7D1A] = 8'h44;
mem[16'h7D1B] = 8'h03;
mem[16'h7D1C] = 8'h0C;
mem[16'h7D1D] = 8'h00;
mem[16'h7D1E] = 8'h44;
mem[16'h7D1F] = 8'h03;
mem[16'h7D20] = 8'h0C;
mem[16'h7D21] = 8'h00;
mem[16'h7D22] = 8'h30;
mem[16'h7D23] = 8'h00;
mem[16'h7D24] = 8'h03;
mem[16'h7D25] = 8'h00;
mem[16'h7D26] = 8'h00;
mem[16'h7D27] = 8'h23;
mem[16'h7D28] = 8'h02;
mem[16'h7D29] = 8'h00;
mem[16'h7D2A] = 8'h00;
mem[16'h7D2B] = 8'h45;
mem[16'h7D2C] = 8'h0A;
mem[16'h7D2D] = 8'h00;
mem[16'h7D2E] = 8'h00;
mem[16'h7D2F] = 8'h15;
mem[16'h7D30] = 8'h00;
mem[16'h7D31] = 8'h00;
mem[16'h7D32] = 8'h40;
mem[16'h7D33] = 8'h0A;
mem[16'h7D34] = 8'h00;
mem[16'h7D35] = 8'h00;
mem[16'h7D36] = 8'h40;
mem[16'h7D37] = 8'h22;
mem[16'h7D38] = 8'h05;
mem[16'h7D39] = 8'h00;
mem[16'h7D3A] = 8'h40;
mem[16'h7D3B] = 8'h11;
mem[16'h7D3C] = 8'h01;
mem[16'h7D3D] = 8'h00;
mem[16'h7D3E] = 8'h18;
mem[16'h7D3F] = 8'h40;
mem[16'h7D40] = 8'h01;
mem[16'h7D41] = 8'h00;
mem[16'h7D42] = 8'h62;
mem[16'h7D43] = 8'h01;
mem[16'h7D44] = 8'h06;
mem[16'h7D45] = 8'h00;
mem[16'h7D46] = 8'h62;
mem[16'h7D47] = 8'h01;
mem[16'h7D48] = 8'h06;
mem[16'h7D49] = 8'h00;
mem[16'h7D4A] = 8'h62;
mem[16'h7D4B] = 8'h01;
mem[16'h7D4C] = 8'h06;
mem[16'h7D4D] = 8'h00;
mem[16'h7D4E] = 8'h18;
mem[16'h7D4F] = 8'h40;
mem[16'h7D50] = 8'h01;
mem[16'h7D51] = 8'h00;
mem[16'h7D52] = 8'h40;
mem[16'h7D53] = 8'h11;
mem[16'h7D54] = 8'h01;
mem[16'h7D55] = 8'h00;
mem[16'h7D56] = 8'h40;
mem[16'h7D57] = 8'h22;
mem[16'h7D58] = 8'h05;
mem[16'h7D59] = 8'h00;
mem[16'h7D5A] = 8'h40;
mem[16'h7D5B] = 8'h0A;
mem[16'h7D5C] = 8'h00;
mem[16'h7D5D] = 8'h00;
mem[16'h7D5E] = 8'h20;
mem[16'h7D5F] = 8'h05;
mem[16'h7D60] = 8'h00;
mem[16'h7D61] = 8'h00;
mem[16'h7D62] = 8'h20;
mem[16'h7D63] = 8'h51;
mem[16'h7D64] = 8'h02;
mem[16'h7D65] = 8'h00;
mem[16'h7D66] = 8'h60;
mem[16'h7D67] = 8'h48;
mem[16'h7D68] = 8'h00;
mem[16'h7D69] = 8'h00;
mem[16'h7D6A] = 8'h0C;
mem[16'h7D6B] = 8'h60;
mem[16'h7D6C] = 8'h00;
mem[16'h7D6D] = 8'h00;
mem[16'h7D6E] = 8'h71;
mem[16'h7D6F] = 8'h00;
mem[16'h7D70] = 8'h03;
mem[16'h7D71] = 8'h00;
mem[16'h7D72] = 8'h71;
mem[16'h7D73] = 8'h00;
mem[16'h7D74] = 8'h03;
mem[16'h7D75] = 8'h00;
mem[16'h7D76] = 8'h71;
mem[16'h7D77] = 8'h00;
mem[16'h7D78] = 8'h03;
mem[16'h7D79] = 8'h00;
mem[16'h7D7A] = 8'h0C;
mem[16'h7D7B] = 8'h60;
mem[16'h7D7C] = 8'h00;
mem[16'h7D7D] = 8'h00;
mem[16'h7D7E] = 8'h60;
mem[16'h7D7F] = 8'h48;
mem[16'h7D80] = 8'h00;
mem[16'h7D81] = 8'h00;
mem[16'h7D82] = 8'h20;
mem[16'h7D83] = 8'h51;
mem[16'h7D84] = 8'h02;
mem[16'h7D85] = 8'h00;
mem[16'h7D86] = 8'h20;
mem[16'h7D87] = 8'h05;
mem[16'h7D88] = 8'h00;
mem[16'h7D89] = 8'h00;
mem[16'h7D8A] = 8'h00;
mem[16'h7D8B] = 8'h50;
mem[16'h7D8C] = 8'h00;
mem[16'h7D8D] = 8'h00;
mem[16'h7D8E] = 8'h00;
mem[16'h7D8F] = 8'h50;
mem[16'h7D90] = 8'h28;
mem[16'h7D91] = 8'h00;
mem[16'h7D92] = 8'h00;
mem[16'h7D93] = 8'h30;
mem[16'h7D94] = 8'h24;
mem[16'h7D95] = 8'h00;
mem[16'h7D96] = 8'h00;
mem[16'h7D97] = 8'h06;
mem[16'h7D98] = 8'h30;
mem[16'h7D99] = 8'h00;
mem[16'h7D9A] = 8'h40;
mem[16'h7D9B] = 8'h38;
mem[16'h7D9C] = 8'h40;
mem[16'h7D9D] = 8'h01;
mem[16'h7D9E] = 8'h40;
mem[16'h7D9F] = 8'h38;
mem[16'h7DA0] = 8'h40;
mem[16'h7DA1] = 8'h01;
mem[16'h7DA2] = 8'h40;
mem[16'h7DA3] = 8'h38;
mem[16'h7DA4] = 8'h40;
mem[16'h7DA5] = 8'h01;
mem[16'h7DA6] = 8'h00;
mem[16'h7DA7] = 8'h06;
mem[16'h7DA8] = 8'h30;
mem[16'h7DA9] = 8'h00;
mem[16'h7DAA] = 8'h00;
mem[16'h7DAB] = 8'h30;
mem[16'h7DAC] = 8'h24;
mem[16'h7DAD] = 8'h00;
mem[16'h7DAE] = 8'h00;
mem[16'h7DAF] = 8'h50;
mem[16'h7DB0] = 8'h28;
mem[16'h7DB1] = 8'h00;
mem[16'h7DB2] = 8'h00;
mem[16'h7DB3] = 8'h50;
mem[16'h7DB4] = 8'h00;
mem[16'h7DB5] = 8'h00;
mem[16'h7DB6] = 8'h00;
mem[16'h7DB7] = 8'h28;
mem[16'h7DB8] = 8'h00;
mem[16'h7DB9] = 8'h00;
mem[16'h7DBA] = 8'h00;
mem[16'h7DBB] = 8'h28;
mem[16'h7DBC] = 8'h14;
mem[16'h7DBD] = 8'h00;
mem[16'h7DBE] = 8'h00;
mem[16'h7DBF] = 8'h18;
mem[16'h7DC0] = 8'h12;
mem[16'h7DC1] = 8'h00;
mem[16'h7DC2] = 8'h00;
mem[16'h7DC3] = 8'h03;
mem[16'h7DC4] = 8'h18;
mem[16'h7DC5] = 8'h00;
mem[16'h7DC6] = 8'h20;
mem[16'h7DC7] = 8'h1C;
mem[16'h7DC8] = 8'h60;
mem[16'h7DC9] = 8'h00;
mem[16'h7DCA] = 8'h20;
mem[16'h7DCB] = 8'h1C;
mem[16'h7DCC] = 8'h60;
mem[16'h7DCD] = 8'h00;
mem[16'h7DCE] = 8'h20;
mem[16'h7DCF] = 8'h1C;
mem[16'h7DD0] = 8'h60;
mem[16'h7DD1] = 8'h00;
mem[16'h7DD2] = 8'h00;
mem[16'h7DD3] = 8'h03;
mem[16'h7DD4] = 8'h18;
mem[16'h7DD5] = 8'h00;
mem[16'h7DD6] = 8'h00;
mem[16'h7DD7] = 8'h18;
mem[16'h7DD8] = 8'h12;
mem[16'h7DD9] = 8'h00;
mem[16'h7DDA] = 8'h00;
mem[16'h7DDB] = 8'h28;
mem[16'h7DDC] = 8'h14;
mem[16'h7DDD] = 8'h00;
mem[16'h7DDE] = 8'h00;
mem[16'h7DDF] = 8'h28;
mem[16'h7DE0] = 8'h00;
mem[16'h7DE1] = 8'h00;
mem[16'h7DE2] = 8'h00;
mem[16'h7DE3] = 8'h14;
mem[16'h7DE4] = 8'h00;
mem[16'h7DE5] = 8'h00;
mem[16'h7DE6] = 8'h00;
mem[16'h7DE7] = 8'h14;
mem[16'h7DE8] = 8'h0A;
mem[16'h7DE9] = 8'h00;
mem[16'h7DEA] = 8'h00;
mem[16'h7DEB] = 8'h0C;
mem[16'h7DEC] = 8'h09;
mem[16'h7DED] = 8'h00;
mem[16'h7DEE] = 8'h40;
mem[16'h7DEF] = 8'h01;
mem[16'h7DF0] = 8'h0C;
mem[16'h7DF1] = 8'h00;
mem[16'h7DF2] = 8'h10;
mem[16'h7DF3] = 8'h0E;
mem[16'h7DF4] = 8'h30;
mem[16'h7DF5] = 8'h00;
mem[16'h7DF6] = 8'h10;
mem[16'h7DF7] = 8'h0E;
mem[16'h7DF8] = 8'h30;
mem[16'h7DF9] = 8'h00;
mem[16'h7DFA] = 8'h10;
mem[16'h7DFB] = 8'h0E;
mem[16'h7DFC] = 8'h30;
mem[16'h7DFD] = 8'h00;
mem[16'h7DFE] = 8'h40;
mem[16'h7DFF] = 8'h01;
mem[16'h7E00] = 8'h0C;
mem[16'h7E01] = 8'h00;
mem[16'h7E02] = 8'h00;
mem[16'h7E03] = 8'h0C;
mem[16'h7E04] = 8'h09;
mem[16'h7E05] = 8'h00;
mem[16'h7E06] = 8'h00;
mem[16'h7E07] = 8'h14;
mem[16'h7E08] = 8'h0A;
mem[16'h7E09] = 8'h00;
mem[16'h7E0A] = 8'h00;
mem[16'h7E0B] = 8'h14;
mem[16'h7E0C] = 8'h00;
mem[16'h7E0D] = 8'h00;
mem[16'h7E0E] = 8'h00;
mem[16'h7E0F] = 8'h0A;
mem[16'h7E10] = 8'h00;
mem[16'h7E11] = 8'h00;
mem[16'h7E12] = 8'h00;
mem[16'h7E13] = 8'h0A;
mem[16'h7E14] = 8'h05;
mem[16'h7E15] = 8'h00;
mem[16'h7E16] = 8'h00;
mem[16'h7E17] = 8'h46;
mem[16'h7E18] = 8'h04;
mem[16'h7E19] = 8'h00;
mem[16'h7E1A] = 8'h60;
mem[16'h7E1B] = 8'h00;
mem[16'h7E1C] = 8'h06;
mem[16'h7E1D] = 8'h00;
mem[16'h7E1E] = 8'h08;
mem[16'h7E1F] = 8'h07;
mem[16'h7E20] = 8'h18;
mem[16'h7E21] = 8'h00;
mem[16'h7E22] = 8'h08;
mem[16'h7E23] = 8'h07;
mem[16'h7E24] = 8'h18;
mem[16'h7E25] = 8'h00;
mem[16'h7E26] = 8'h08;
mem[16'h7E27] = 8'h07;
mem[16'h7E28] = 8'h18;
mem[16'h7E29] = 8'h00;
mem[16'h7E2A] = 8'h60;
mem[16'h7E2B] = 8'h00;
mem[16'h7E2C] = 8'h06;
mem[16'h7E2D] = 8'h00;
mem[16'h7E2E] = 8'h00;
mem[16'h7E2F] = 8'h46;
mem[16'h7E30] = 8'h04;
mem[16'h7E31] = 8'h00;
mem[16'h7E32] = 8'h00;
mem[16'h7E33] = 8'h0A;
mem[16'h7E34] = 8'h05;
mem[16'h7E35] = 8'h00;
mem[16'h7E36] = 8'h00;
mem[16'h7E37] = 8'h0A;
mem[16'h7E38] = 8'h00;
mem[16'h7E39] = 8'h00;
mem[16'h7E3A] = 8'h00;
mem[16'h7E3B] = 8'h05;
mem[16'h7E3C] = 8'h00;
mem[16'h7E3D] = 8'h00;
mem[16'h7E3E] = 8'h00;
mem[16'h7E3F] = 8'h45;
mem[16'h7E40] = 8'h02;
mem[16'h7E41] = 8'h00;
mem[16'h7E42] = 8'h00;
mem[16'h7E43] = 8'h23;
mem[16'h7E44] = 8'h02;
mem[16'h7E45] = 8'h00;
mem[16'h7E46] = 8'h30;
mem[16'h7E47] = 8'h00;
mem[16'h7E48] = 8'h03;
mem[16'h7E49] = 8'h00;
mem[16'h7E4A] = 8'h44;
mem[16'h7E4B] = 8'h03;
mem[16'h7E4C] = 8'h0C;
mem[16'h7E4D] = 8'h00;
mem[16'h7E4E] = 8'h44;
mem[16'h7E4F] = 8'h03;
mem[16'h7E50] = 8'h0C;
mem[16'h7E51] = 8'h00;
mem[16'h7E52] = 8'h44;
mem[16'h7E53] = 8'h03;
mem[16'h7E54] = 8'h0C;
mem[16'h7E55] = 8'h00;
mem[16'h7E56] = 8'h30;
mem[16'h7E57] = 8'h00;
mem[16'h7E58] = 8'h03;
mem[16'h7E59] = 8'h00;
mem[16'h7E5A] = 8'h00;
mem[16'h7E5B] = 8'h23;
mem[16'h7E5C] = 8'h02;
mem[16'h7E5D] = 8'h00;
mem[16'h7E5E] = 8'h00;
mem[16'h7E5F] = 8'h45;
mem[16'h7E60] = 8'h02;
mem[16'h7E61] = 8'h00;
mem[16'h7E62] = 8'h00;
mem[16'h7E63] = 8'h05;
mem[16'h7E64] = 8'h00;
mem[16'h7E65] = 8'h00;
mem[16'h7E66] = 8'h40;
mem[16'h7E67] = 8'h02;
mem[16'h7E68] = 8'h00;
mem[16'h7E69] = 8'h00;
mem[16'h7E6A] = 8'h40;
mem[16'h7E6B] = 8'h22;
mem[16'h7E6C] = 8'h01;
mem[16'h7E6D] = 8'h00;
mem[16'h7E6E] = 8'h40;
mem[16'h7E6F] = 8'h11;
mem[16'h7E70] = 8'h01;
mem[16'h7E71] = 8'h00;
mem[16'h7E72] = 8'h18;
mem[16'h7E73] = 8'h40;
mem[16'h7E74] = 8'h01;
mem[16'h7E75] = 8'h00;
mem[16'h7E76] = 8'h62;
mem[16'h7E77] = 8'h01;
mem[16'h7E78] = 8'h06;
mem[16'h7E79] = 8'h00;
mem[16'h7E7A] = 8'h62;
mem[16'h7E7B] = 8'h01;
mem[16'h7E7C] = 8'h06;
mem[16'h7E7D] = 8'h00;
mem[16'h7E7E] = 8'h62;
mem[16'h7E7F] = 8'h01;
mem[16'h7E80] = 8'h06;
mem[16'h7E81] = 8'h00;
mem[16'h7E82] = 8'h18;
mem[16'h7E83] = 8'h40;
mem[16'h7E84] = 8'h01;
mem[16'h7E85] = 8'h00;
mem[16'h7E86] = 8'h40;
mem[16'h7E87] = 8'h11;
mem[16'h7E88] = 8'h01;
mem[16'h7E89] = 8'h00;
mem[16'h7E8A] = 8'h40;
mem[16'h7E8B] = 8'h22;
mem[16'h7E8C] = 8'h01;
mem[16'h7E8D] = 8'h00;
mem[16'h7E8E] = 8'h40;
mem[16'h7E8F] = 8'h02;
mem[16'h7E90] = 8'h00;
mem[16'h7E91] = 8'h00;
mem[16'h7E92] = 8'h20;
mem[16'h7E93] = 8'h01;
mem[16'h7E94] = 8'h00;
mem[16'h7E95] = 8'h00;
mem[16'h7E96] = 8'h20;
mem[16'h7E97] = 8'h51;
mem[16'h7E98] = 8'h00;
mem[16'h7E99] = 8'h00;
mem[16'h7E9A] = 8'h60;
mem[16'h7E9B] = 8'h48;
mem[16'h7E9C] = 8'h00;
mem[16'h7E9D] = 8'h00;
mem[16'h7E9E] = 8'h0C;
mem[16'h7E9F] = 8'h60;
mem[16'h7EA0] = 8'h00;
mem[16'h7EA1] = 8'h00;
mem[16'h7EA2] = 8'h71;
mem[16'h7EA3] = 8'h00;
mem[16'h7EA4] = 8'h03;
mem[16'h7EA5] = 8'h00;
mem[16'h7EA6] = 8'h71;
mem[16'h7EA7] = 8'h00;
mem[16'h7EA8] = 8'h03;
mem[16'h7EA9] = 8'h00;
mem[16'h7EAA] = 8'h71;
mem[16'h7EAB] = 8'h00;
mem[16'h7EAC] = 8'h03;
mem[16'h7EAD] = 8'h00;
mem[16'h7EAE] = 8'h0C;
mem[16'h7EAF] = 8'h60;
mem[16'h7EB0] = 8'h00;
mem[16'h7EB1] = 8'h00;
mem[16'h7EB2] = 8'h60;
mem[16'h7EB3] = 8'h48;
mem[16'h7EB4] = 8'h00;
mem[16'h7EB5] = 8'h00;
mem[16'h7EB6] = 8'h20;
mem[16'h7EB7] = 8'h51;
mem[16'h7EB8] = 8'h00;
mem[16'h7EB9] = 8'h00;
mem[16'h7EBA] = 8'h20;
mem[16'h7EBB] = 8'h01;
mem[16'h7EBC] = 8'h00;
mem[16'h7EBD] = 8'h00;
mem[16'h7EBE] = 8'hA9;
mem[16'h7EBF] = 8'hDB;
mem[16'h7EC0] = 8'hA0;
mem[16'h7EC1] = 8'h7E;
mem[16'h7EC2] = 8'h20;
mem[16'h7EC3] = 8'h42;
mem[16'h7EC4] = 8'h6A;
mem[16'h7EC5] = 8'hA9;
mem[16'h7EC6] = 8'h26;
mem[16'h7EC7] = 8'h8D;
mem[16'h7EC8] = 8'hF9;
mem[16'h7EC9] = 8'h69;
mem[16'h7ECA] = 8'hAD;
mem[16'h7ECB] = 8'hCF;
mem[16'h7ECC] = 8'h4D;
mem[16'h7ECD] = 8'h85;
mem[16'h7ECE] = 8'h57;
mem[16'h7ECF] = 8'hAD;
mem[16'h7ED0] = 8'hD0;
mem[16'h7ED1] = 8'h4D;
mem[16'h7ED2] = 8'h38;
mem[16'h7ED3] = 8'hE9;
mem[16'h7ED4] = 8'h03;
mem[16'h7ED5] = 8'h85;
mem[16'h7ED6] = 8'h56;
mem[16'h7ED7] = 8'h20;
mem[16'h7ED8] = 8'h33;
mem[16'h7ED9] = 8'h69;
mem[16'h7EDA] = 8'h60;
mem[16'h7EDB] = 8'h00;
mem[16'h7EDC] = 8'h00;
mem[16'h7EDD] = 8'h60;
mem[16'h7EDE] = 8'h03;
mem[16'h7EDF] = 8'h70;
mem[16'h7EE0] = 8'h07;
mem[16'h7EE1] = 8'h48;
mem[16'h7EE2] = 8'h09;
mem[16'h7EE3] = 8'h48;
mem[16'h7EE4] = 8'h09;
mem[16'h7EE5] = 8'h78;
mem[16'h7EE6] = 8'h0F;
mem[16'h7EE7] = 8'h78;
mem[16'h7EE8] = 8'h0F;
mem[16'h7EE9] = 8'h33;
mem[16'h7EEA] = 8'h66;
mem[16'h7EEB] = 8'h33;
mem[16'h7EEC] = 8'h66;
mem[16'h7EED] = 8'h72;
mem[16'h7EEE] = 8'h27;
mem[16'h7EEF] = 8'h24;
mem[16'h7EF0] = 8'h12;
mem[16'h7EF1] = 8'h48;
mem[16'h7EF2] = 8'h09;
mem[16'h7EF3] = 8'h10;
mem[16'h7EF4] = 8'h04;
mem[16'h7EF5] = 8'h20;
mem[16'h7EF6] = 8'h02;
mem[16'h7EF7] = 8'h40;
mem[16'h7EF8] = 8'h01;
mem[16'h7EF9] = 8'h40;
mem[16'h7EFA] = 8'h01;
mem[16'h7EFB] = 8'h20;
mem[16'h7EFC] = 8'h02;
mem[16'h7EFD] = 8'h18;
mem[16'h7EFE] = 8'h0C;
mem[16'h7EFF] = 8'h18;
mem[16'h7F00] = 8'h0C;
mem[16'h7F01] = 8'hAD;
mem[16'h7F02] = 8'h00;
mem[16'h7F03] = 8'hC0;
mem[16'h7F04] = 8'hC9;
mem[16'h7F05] = 8'hA1;
mem[16'h7F06] = 8'hD0;
mem[16'h7F07] = 8'h35;
mem[16'h7F08] = 8'hAD;
mem[16'h7F09] = 8'h4F;
mem[16'h7F0A] = 8'h7F;
mem[16'h7F0B] = 8'h49;
mem[16'h7F0C] = 8'h01;
mem[16'h7F0D] = 8'h8D;
mem[16'h7F0E] = 8'h4F;
mem[16'h7F0F] = 8'h7F;
mem[16'h7F10] = 8'h0A;
mem[16'h7F11] = 8'h18;
mem[16'h7F12] = 8'h69;
mem[16'h7F13] = 8'h06;
mem[16'h7F14] = 8'h8D;
mem[16'h7F15] = 8'hE0;
mem[16'h7F16] = 8'h91;
mem[16'h7F17] = 8'hA9;
mem[16'h7F18] = 8'h17;
mem[16'h7F19] = 8'h85;
mem[16'h7F1A] = 8'h25;
mem[16'h7F1B] = 8'hA9;
mem[16'h7F1C] = 8'h25;
mem[16'h7F1D] = 8'h85;
mem[16'h7F1E] = 8'h24;
mem[16'h7F1F] = 8'hAD;
mem[16'h7F20] = 8'h50;
mem[16'h7F21] = 8'h7F;
mem[16'h7F22] = 8'h20;
mem[16'h7F23] = 8'hED;
mem[16'h7F24] = 8'hFD;
mem[16'h7F25] = 8'hC6;
mem[16'h7F26] = 8'h24;
mem[16'h7F27] = 8'hAD;
mem[16'h7F28] = 8'h51;
mem[16'h7F29] = 8'h7F;
mem[16'h7F2A] = 8'h85;
mem[16'h7F2B] = 8'h60;
mem[16'h7F2C] = 8'h20;
mem[16'h7F2D] = 8'hED;
mem[16'h7F2E] = 8'hFD;
mem[16'h7F2F] = 8'hAD;
mem[16'h7F30] = 8'h50;
mem[16'h7F31] = 8'h7F;
mem[16'h7F32] = 8'h8D;
mem[16'h7F33] = 8'h51;
mem[16'h7F34] = 8'h7F;
mem[16'h7F35] = 8'hA5;
mem[16'h7F36] = 8'h60;
mem[16'h7F37] = 8'h8D;
mem[16'h7F38] = 8'h50;
mem[16'h7F39] = 8'h7F;
mem[16'h7F3A] = 8'hAD;
mem[16'h7F3B] = 8'h10;
mem[16'h7F3C] = 8'hC0;
mem[16'h7F3D] = 8'hAD;
mem[16'h7F3E] = 8'h4F;
mem[16'h7F3F] = 8'h7F;
mem[16'h7F40] = 8'hD0;
mem[16'h7F41] = 8'h01;
mem[16'h7F42] = 8'h60;
mem[16'h7F43] = 8'hA9;
mem[16'h7F44] = 8'h78;
mem[16'h7F45] = 8'h20;
mem[16'h7F46] = 8'hA8;
mem[16'h7F47] = 8'hFC;
mem[16'h7F48] = 8'h20;
mem[16'h7F49] = 8'hBD;
mem[16'h7F4A] = 8'h4A;
mem[16'h7F4B] = 8'h20;
mem[16'h7F4C] = 8'hD4;
mem[16'h7F4D] = 8'h90;
mem[16'h7F4E] = 8'h60;
mem[16'h7F4F] = 8'h00;
mem[16'h7F50] = 8'hCE;
mem[16'h7F51] = 8'hD3;
mem[16'h7F52] = 8'hA2;
mem[16'h7F53] = 8'h01;
mem[16'h7F54] = 8'h20;
mem[16'h7F55] = 8'h1E;
mem[16'h7F56] = 8'hFB;
mem[16'h7F57] = 8'hAD;
mem[16'h7F58] = 8'hCD;
mem[16'h7F59] = 8'h7F;
mem[16'h7F5A] = 8'hC5;
mem[16'h7F5B] = 8'h89;
mem[16'h7F5C] = 8'h90;
mem[16'h7F5D] = 8'h11;
mem[16'h7F5E] = 8'hC5;
mem[16'h7F5F] = 8'h8A;
mem[16'h7F60] = 8'hB0;
mem[16'h7F61] = 8'h0D;
mem[16'h7F62] = 8'hC4;
mem[16'h7F63] = 8'h89;
mem[16'h7F64] = 8'h90;
mem[16'h7F65] = 8'h09;
mem[16'h7F66] = 8'hC4;
mem[16'h7F67] = 8'h8A;
mem[16'h7F68] = 8'hB0;
mem[16'h7F69] = 8'h05;
mem[16'h7F6A] = 8'hA9;
mem[16'h7F6B] = 8'h00;
mem[16'h7F6C] = 8'h85;
mem[16'h7F6D] = 8'h86;
mem[16'h7F6E] = 8'h60;
mem[16'h7F6F] = 8'hA6;
mem[16'h7F70] = 8'h86;
mem[16'h7F71] = 8'hD0;
mem[16'h7F72] = 8'hFB;
mem[16'h7F73] = 8'h38;
mem[16'h7F74] = 8'hE9;
mem[16'h7F75] = 8'h80;
mem[16'h7F76] = 8'h8D;
mem[16'h7F77] = 8'hCE;
mem[16'h7F78] = 8'h7F;
mem[16'h7F79] = 8'h98;
mem[16'h7F7A] = 8'h49;
mem[16'h7F7B] = 8'hFF;
mem[16'h7F7C] = 8'h38;
mem[16'h7F7D] = 8'hE9;
mem[16'h7F7E] = 8'h80;
mem[16'h7F7F] = 8'h8D;
mem[16'h7F80] = 8'hCF;
mem[16'h7F81] = 8'h7F;
mem[16'h7F82] = 8'h10;
mem[16'h7F83] = 8'h2C;
mem[16'h7F84] = 8'hAD;
mem[16'h7F85] = 8'hCE;
mem[16'h7F86] = 8'h7F;
mem[16'h7F87] = 8'h30;
mem[16'h7F88] = 8'h18;
mem[16'h7F89] = 8'h18;
mem[16'h7F8A] = 8'h6D;
mem[16'h7F8B] = 8'hCF;
mem[16'h7F8C] = 8'h7F;
mem[16'h7F8D] = 8'h10;
mem[16'h7F8E] = 8'h09;
mem[16'h7F8F] = 8'h68;
mem[16'h7F90] = 8'h68;
mem[16'h7F91] = 8'hA5;
mem[16'h7F92] = 8'h7E;
mem[16'h7F93] = 8'h85;
mem[16'h7F94] = 8'h86;
mem[16'h7F95] = 8'h4C;
mem[16'h7F96] = 8'hF2;
mem[16'h7F97] = 8'h4A;
mem[16'h7F98] = 8'h68;
mem[16'h7F99] = 8'h68;
mem[16'h7F9A] = 8'hA5;
mem[16'h7F9B] = 8'h80;
mem[16'h7F9C] = 8'h85;
mem[16'h7F9D] = 8'h86;
mem[16'h7F9E] = 8'h4C;
mem[16'h7F9F] = 8'h39;
mem[16'h7FA0] = 8'h4B;
mem[16'h7FA1] = 8'h38;
mem[16'h7FA2] = 8'hED;
mem[16'h7FA3] = 8'hCF;
mem[16'h7FA4] = 8'h7F;
mem[16'h7FA5] = 8'h10;
mem[16'h7FA6] = 8'hE8;
mem[16'h7FA7] = 8'h68;
mem[16'h7FA8] = 8'h68;
mem[16'h7FA9] = 8'hA5;
mem[16'h7FAA] = 8'h7F;
mem[16'h7FAB] = 8'h85;
mem[16'h7FAC] = 8'h86;
mem[16'h7FAD] = 8'h4C;
mem[16'h7FAE] = 8'h19;
mem[16'h7FAF] = 8'h4B;
mem[16'h7FB0] = 8'hAD;
mem[16'h7FB1] = 8'hCE;
mem[16'h7FB2] = 8'h7F;
mem[16'h7FB3] = 8'h30;
mem[16'h7FB4] = 8'h0F;
mem[16'h7FB5] = 8'h38;
mem[16'h7FB6] = 8'hED;
mem[16'h7FB7] = 8'hCF;
mem[16'h7FB8] = 8'h7F;
mem[16'h7FB9] = 8'h10;
mem[16'h7FBA] = 8'hDD;
mem[16'h7FBB] = 8'h68;
mem[16'h7FBC] = 8'h68;
mem[16'h7FBD] = 8'hA5;
mem[16'h7FBE] = 8'h7D;
mem[16'h7FBF] = 8'h85;
mem[16'h7FC0] = 8'h86;
mem[16'h7FC1] = 8'h4C;
mem[16'h7FC2] = 8'hD2;
mem[16'h7FC3] = 8'h4A;
mem[16'h7FC4] = 8'h18;
mem[16'h7FC5] = 8'h6D;
mem[16'h7FC6] = 8'hCF;
mem[16'h7FC7] = 8'h7F;
mem[16'h7FC8] = 8'h10;
mem[16'h7FC9] = 8'hF1;
mem[16'h7FCA] = 8'h4C;
mem[16'h7FCB] = 8'hA7;
mem[16'h7FCC] = 8'h7F;
mem[16'h7FCD] = 8'h00;
mem[16'h7FCE] = 8'h00;
mem[16'h7FCF] = 8'h00;
mem[16'h7FD0] = 8'hA5;
mem[16'h7FD1] = 8'h85;
mem[16'h7FD2] = 8'hF0;
mem[16'h7FD3] = 8'h08;
mem[16'h7FD4] = 8'hA2;
mem[16'h7FD5] = 8'h00;
mem[16'h7FD6] = 8'h20;
mem[16'h7FD7] = 8'h1E;
mem[16'h7FD8] = 8'hFB;
mem[16'h7FD9] = 8'h8C;
mem[16'h7FDA] = 8'hCD;
mem[16'h7FDB] = 8'h7F;
mem[16'h7FDC] = 8'h60;
mem[16'h7FDD] = 8'h31;
mem[16'h7FDE] = 8'h37;
mem[16'h7FDF] = 8'h31;
mem[16'h7FE0] = 8'h45;
mem[16'h7FE1] = 8'h35;
mem[16'h7FE2] = 8'h38;
mem[16'h7FE3] = 8'h31;
mem[16'h7FE4] = 8'h37;
mem[16'h7FE5] = 8'h33;
mem[16'h7FE6] = 8'h30;
mem[16'h7FE7] = 8'h0D;
mem[16'h7FE8] = 8'h17;
mem[16'h7FE9] = 8'hE4;
mem[16'h7FEA] = 8'h20;
mem[16'h7FEB] = 8'h31;
mem[16'h7FEC] = 8'h37;
mem[16'h7FED] = 8'h33;
mem[16'h7FEE] = 8'h30;
mem[16'h7FEF] = 8'h31;
mem[16'h7FF0] = 8'h37;
mem[16'h7FF1] = 8'h33;
mem[16'h7FF2] = 8'h30;
mem[16'h7FF3] = 8'h31;
mem[16'h7FF4] = 8'h45;
mem[16'h7FF5] = 8'h35;
mem[16'h7FF6] = 8'h38;
mem[16'h7FF7] = 8'h36;
mem[16'h7FF8] = 8'h30;
mem[16'h7FF9] = 8'h31;
mem[16'h7FFA] = 8'h37;
mem[16'h7FFB] = 8'h32;
mem[16'h7FFC] = 8'h38;
mem[16'h7FFD] = 8'h34;
mem[16'h7FFE] = 8'h30;
mem[16'h7FFF] = 8'h0D;
mem[16'h8000] = 8'h40;
mem[16'h8001] = 8'h00;
mem[16'h8002] = 8'h00;
mem[16'h8003] = 8'h40;
mem[16'h8004] = 8'h01;
mem[16'h8005] = 8'h00;
mem[16'h8006] = 8'h41;
mem[16'h8007] = 8'h02;
mem[16'h8008] = 8'h01;
mem[16'h8009] = 8'h45;
mem[16'h800A] = 8'h02;
mem[16'h800B] = 8'h01;
mem[16'h800C] = 8'h54;
mem[16'h800D] = 8'h22;
mem[16'h800E] = 8'h00;
mem[16'h800F] = 8'h54;
mem[16'h8010] = 8'h2A;
mem[16'h8011] = 8'h00;
mem[16'h8012] = 8'h50;
mem[16'h8013] = 8'h2A;
mem[16'h8014] = 8'h00;
mem[16'h8015] = 8'h50;
mem[16'h8016] = 8'h2A;
mem[16'h8017] = 8'h00;
mem[16'h8018] = 8'h50;
mem[16'h8019] = 8'h0A;
mem[16'h801A] = 8'h00;
mem[16'h801B] = 8'h55;
mem[16'h801C] = 8'h0A;
mem[16'h801D] = 8'h00;
mem[16'h801E] = 8'h55;
mem[16'h801F] = 8'h2A;
mem[16'h8020] = 8'h00;
mem[16'h8021] = 8'h50;
mem[16'h8022] = 8'h2A;
mem[16'h8023] = 8'h01;
mem[16'h8024] = 8'h40;
mem[16'h8025] = 8'h2A;
mem[16'h8026] = 8'h05;
mem[16'h8027] = 8'h40;
mem[16'h8028] = 8'h02;
mem[16'h8029] = 8'h05;
mem[16'h802A] = 8'h40;
mem[16'h802B] = 8'h02;
mem[16'h802C] = 8'h00;
mem[16'h802D] = 8'h00;
mem[16'h802E] = 8'h03;
mem[16'h802F] = 8'h00;
mem[16'h8030] = 8'h00;
mem[16'h8031] = 8'h02;
mem[16'h8032] = 8'h00;
mem[16'h8033] = 8'h06;
mem[16'h8034] = 8'h00;
mem[16'h8035] = 8'h18;
mem[16'h8036] = 8'h00;
mem[16'h8037] = 8'h60;
mem[16'h8038] = 8'h00;
mem[16'h8039] = 8'h60;
mem[16'h803A] = 8'h00;
mem[16'h803B] = 8'h60;
mem[16'h803C] = 8'h00;
mem[16'h803D] = 8'h60;
mem[16'h803E] = 8'h00;
mem[16'h803F] = 8'h60;
mem[16'h8040] = 8'h00;
mem[16'h8041] = 8'h18;
mem[16'h8042] = 8'h00;
mem[16'h8043] = 8'h06;
mem[16'h8044] = 8'h00;
mem[16'h8045] = 8'h0C;
mem[16'h8046] = 8'h00;
mem[16'h8047] = 8'h30;
mem[16'h8048] = 8'h00;
mem[16'h8049] = 8'h40;
mem[16'h804A] = 8'h01;
mem[16'h804B] = 8'h40;
mem[16'h804C] = 8'h01;
mem[16'h804D] = 8'h40;
mem[16'h804E] = 8'h01;
mem[16'h804F] = 8'h40;
mem[16'h8050] = 8'h01;
mem[16'h8051] = 8'h40;
mem[16'h8052] = 8'h01;
mem[16'h8053] = 8'h30;
mem[16'h8054] = 8'h00;
mem[16'h8055] = 8'h0C;
mem[16'h8056] = 8'h00;
mem[16'h8057] = 8'h18;
mem[16'h8058] = 8'h00;
mem[16'h8059] = 8'h60;
mem[16'h805A] = 8'h00;
mem[16'h805B] = 8'h00;
mem[16'h805C] = 8'h03;
mem[16'h805D] = 8'h00;
mem[16'h805E] = 8'h03;
mem[16'h805F] = 8'h00;
mem[16'h8060] = 8'h03;
mem[16'h8061] = 8'h00;
mem[16'h8062] = 8'h03;
mem[16'h8063] = 8'h00;
mem[16'h8064] = 8'h03;
mem[16'h8065] = 8'h60;
mem[16'h8066] = 8'h00;
mem[16'h8067] = 8'h18;
mem[16'h8068] = 8'h00;
mem[16'h8069] = 8'h30;
mem[16'h806A] = 8'h00;
mem[16'h806B] = 8'h40;
mem[16'h806C] = 8'h01;
mem[16'h806D] = 8'h00;
mem[16'h806E] = 8'h06;
mem[16'h806F] = 8'h00;
mem[16'h8070] = 8'h06;
mem[16'h8071] = 8'h00;
mem[16'h8072] = 8'h06;
mem[16'h8073] = 8'h00;
mem[16'h8074] = 8'h06;
mem[16'h8075] = 8'h00;
mem[16'h8076] = 8'h06;
mem[16'h8077] = 8'h40;
mem[16'h8078] = 8'h01;
mem[16'h8079] = 8'h30;
mem[16'h807A] = 8'h00;
mem[16'h807B] = 8'h60;
mem[16'h807C] = 8'h00;
mem[16'h807D] = 8'h00;
mem[16'h807E] = 8'h03;
mem[16'h807F] = 8'h00;
mem[16'h8080] = 8'h0C;
mem[16'h8081] = 8'h00;
mem[16'h8082] = 8'h0C;
mem[16'h8083] = 8'h00;
mem[16'h8084] = 8'h0C;
mem[16'h8085] = 8'h00;
mem[16'h8086] = 8'h0C;
mem[16'h8087] = 8'h00;
mem[16'h8088] = 8'h0C;
mem[16'h8089] = 8'h00;
mem[16'h808A] = 8'h03;
mem[16'h808B] = 8'h60;
mem[16'h808C] = 8'h00;
mem[16'h808D] = 8'h40;
mem[16'h808E] = 8'h01;
mem[16'h808F] = 8'h00;
mem[16'h8090] = 8'h06;
mem[16'h8091] = 8'h00;
mem[16'h8092] = 8'h18;
mem[16'h8093] = 8'h00;
mem[16'h8094] = 8'h18;
mem[16'h8095] = 8'h00;
mem[16'h8096] = 8'h18;
mem[16'h8097] = 8'h00;
mem[16'h8098] = 8'h18;
mem[16'h8099] = 8'h00;
mem[16'h809A] = 8'h18;
mem[16'h809B] = 8'h00;
mem[16'h809C] = 8'h06;
mem[16'h809D] = 8'h40;
mem[16'h809E] = 8'h01;
mem[16'h809F] = 8'h00;
mem[16'h80A0] = 8'h03;
mem[16'h80A1] = 8'h00;
mem[16'h80A2] = 8'h0C;
mem[16'h80A3] = 8'h00;
mem[16'h80A4] = 8'h30;
mem[16'h80A5] = 8'h00;
mem[16'h80A6] = 8'h30;
mem[16'h80A7] = 8'h00;
mem[16'h80A8] = 8'h30;
mem[16'h80A9] = 8'h00;
mem[16'h80AA] = 8'h30;
mem[16'h80AB] = 8'h00;
mem[16'h80AC] = 8'h30;
mem[16'h80AD] = 8'h00;
mem[16'h80AE] = 8'h0C;
mem[16'h80AF] = 8'h00;
mem[16'h80B0] = 8'h03;
mem[16'h80B1] = 8'h1E;
mem[16'h80B2] = 8'h00;
mem[16'h80B3] = 8'h00;
mem[16'h80B4] = 8'h78;
mem[16'h80B5] = 8'h00;
mem[16'h80B6] = 8'h00;
mem[16'h80B7] = 8'h60;
mem[16'h80B8] = 8'h03;
mem[16'h80B9] = 8'h00;
mem[16'h80BA] = 8'h60;
mem[16'h80BB] = 8'h03;
mem[16'h80BC] = 8'h00;
mem[16'h80BD] = 8'h60;
mem[16'h80BE] = 8'h03;
mem[16'h80BF] = 8'h00;
mem[16'h80C0] = 8'h60;
mem[16'h80C1] = 8'h03;
mem[16'h80C2] = 8'h00;
mem[16'h80C3] = 8'h60;
mem[16'h80C4] = 8'h03;
mem[16'h80C5] = 8'h00;
mem[16'h80C6] = 8'h78;
mem[16'h80C7] = 8'h00;
mem[16'h80C8] = 8'h00;
mem[16'h80C9] = 8'h1E;
mem[16'h80CA] = 8'h00;
mem[16'h80CB] = 8'h00;
mem[16'h80CC] = 8'h3C;
mem[16'h80CD] = 8'h00;
mem[16'h80CE] = 8'h00;
mem[16'h80CF] = 8'h70;
mem[16'h80D0] = 8'h01;
mem[16'h80D1] = 8'h00;
mem[16'h80D2] = 8'h40;
mem[16'h80D3] = 8'h07;
mem[16'h80D4] = 8'h00;
mem[16'h80D5] = 8'h40;
mem[16'h80D6] = 8'h07;
mem[16'h80D7] = 8'h00;
mem[16'h80D8] = 8'h40;
mem[16'h80D9] = 8'h07;
mem[16'h80DA] = 8'h00;
mem[16'h80DB] = 8'h40;
mem[16'h80DC] = 8'h07;
mem[16'h80DD] = 8'h00;
mem[16'h80DE] = 8'h40;
mem[16'h80DF] = 8'h07;
mem[16'h80E0] = 8'h00;
mem[16'h80E1] = 8'h70;
mem[16'h80E2] = 8'h01;
mem[16'h80E3] = 8'h00;
mem[16'h80E4] = 8'h3C;
mem[16'h80E5] = 8'h00;
mem[16'h80E6] = 8'h00;
mem[16'h80E7] = 8'h78;
mem[16'h80E8] = 8'h00;
mem[16'h80E9] = 8'h00;
mem[16'h80EA] = 8'h60;
mem[16'h80EB] = 8'h03;
mem[16'h80EC] = 8'h00;
mem[16'h80ED] = 8'h00;
mem[16'h80EE] = 8'h0F;
mem[16'h80EF] = 8'h00;
mem[16'h80F0] = 8'h00;
mem[16'h80F1] = 8'h0F;
mem[16'h80F2] = 8'h00;
mem[16'h80F3] = 8'h00;
mem[16'h80F4] = 8'h0F;
mem[16'h80F5] = 8'h00;
mem[16'h80F6] = 8'h00;
mem[16'h80F7] = 8'h0F;
mem[16'h80F8] = 8'h00;
mem[16'h80F9] = 8'h00;
mem[16'h80FA] = 8'h0F;
mem[16'h80FB] = 8'h00;
mem[16'h80FC] = 8'h60;
mem[16'h80FD] = 8'h03;
mem[16'h80FE] = 8'h00;
mem[16'h80FF] = 8'h78;
mem[16'h8100] = 8'h00;
mem[16'h8101] = 8'h00;
mem[16'h8102] = 8'h70;
mem[16'h8103] = 8'h01;
mem[16'h8104] = 8'h00;
mem[16'h8105] = 8'h40;
mem[16'h8106] = 8'h07;
mem[16'h8107] = 8'h00;
mem[16'h8108] = 8'h00;
mem[16'h8109] = 8'h1E;
mem[16'h810A] = 8'h00;
mem[16'h810B] = 8'h00;
mem[16'h810C] = 8'h1E;
mem[16'h810D] = 8'h00;
mem[16'h810E] = 8'h00;
mem[16'h810F] = 8'h1E;
mem[16'h8110] = 8'h00;
mem[16'h8111] = 8'h00;
mem[16'h8112] = 8'h1E;
mem[16'h8113] = 8'h00;
mem[16'h8114] = 8'h00;
mem[16'h8115] = 8'h1E;
mem[16'h8116] = 8'h00;
mem[16'h8117] = 8'h40;
mem[16'h8118] = 8'h07;
mem[16'h8119] = 8'h00;
mem[16'h811A] = 8'h70;
mem[16'h811B] = 8'h01;
mem[16'h811C] = 8'h00;
mem[16'h811D] = 8'h60;
mem[16'h811E] = 8'h03;
mem[16'h811F] = 8'h00;
mem[16'h8120] = 8'h00;
mem[16'h8121] = 8'h0F;
mem[16'h8122] = 8'h00;
mem[16'h8123] = 8'h00;
mem[16'h8124] = 8'h3C;
mem[16'h8125] = 8'h00;
mem[16'h8126] = 8'h00;
mem[16'h8127] = 8'h3C;
mem[16'h8128] = 8'h00;
mem[16'h8129] = 8'h00;
mem[16'h812A] = 8'h3C;
mem[16'h812B] = 8'h00;
mem[16'h812C] = 8'h00;
mem[16'h812D] = 8'h3C;
mem[16'h812E] = 8'h00;
mem[16'h812F] = 8'h00;
mem[16'h8130] = 8'h3C;
mem[16'h8131] = 8'h00;
mem[16'h8132] = 8'h00;
mem[16'h8133] = 8'h0F;
mem[16'h8134] = 8'h00;
mem[16'h8135] = 8'h60;
mem[16'h8136] = 8'h03;
mem[16'h8137] = 8'h00;
mem[16'h8138] = 8'h40;
mem[16'h8139] = 8'h07;
mem[16'h813A] = 8'h00;
mem[16'h813B] = 8'h00;
mem[16'h813C] = 8'h1E;
mem[16'h813D] = 8'h00;
mem[16'h813E] = 8'h00;
mem[16'h813F] = 8'h78;
mem[16'h8140] = 8'h00;
mem[16'h8141] = 8'h00;
mem[16'h8142] = 8'h78;
mem[16'h8143] = 8'h00;
mem[16'h8144] = 8'h00;
mem[16'h8145] = 8'h78;
mem[16'h8146] = 8'h00;
mem[16'h8147] = 8'h00;
mem[16'h8148] = 8'h78;
mem[16'h8149] = 8'h00;
mem[16'h814A] = 8'h00;
mem[16'h814B] = 8'h78;
mem[16'h814C] = 8'h00;
mem[16'h814D] = 8'h00;
mem[16'h814E] = 8'h1E;
mem[16'h814F] = 8'h00;
mem[16'h8150] = 8'h40;
mem[16'h8151] = 8'h07;
mem[16'h8152] = 8'h00;
mem[16'h8153] = 8'h00;
mem[16'h8154] = 8'h0F;
mem[16'h8155] = 8'h00;
mem[16'h8156] = 8'h00;
mem[16'h8157] = 8'h3C;
mem[16'h8158] = 8'h00;
mem[16'h8159] = 8'h00;
mem[16'h815A] = 8'h70;
mem[16'h815B] = 8'h01;
mem[16'h815C] = 8'h00;
mem[16'h815D] = 8'h70;
mem[16'h815E] = 8'h01;
mem[16'h815F] = 8'h00;
mem[16'h8160] = 8'h70;
mem[16'h8161] = 8'h01;
mem[16'h8162] = 8'h00;
mem[16'h8163] = 8'h70;
mem[16'h8164] = 8'h01;
mem[16'h8165] = 8'h00;
mem[16'h8166] = 8'h70;
mem[16'h8167] = 8'h01;
mem[16'h8168] = 8'h00;
mem[16'h8169] = 8'h3C;
mem[16'h816A] = 8'h00;
mem[16'h816B] = 8'h00;
mem[16'h816C] = 8'h0F;
mem[16'h816D] = 8'h00;
mem[16'h816E] = 8'h20;
mem[16'h816F] = 8'h10;
mem[16'h8170] = 8'h00;
mem[16'h8171] = 8'h00;
mem[16'h8172] = 8'h28;
mem[16'h8173] = 8'h50;
mem[16'h8174] = 8'h00;
mem[16'h8175] = 8'h00;
mem[16'h8176] = 8'h00;
mem[16'h8177] = 8'h00;
mem[16'h8178] = 8'h00;
mem[16'h8179] = 8'h00;
mem[16'h817A] = 8'h6A;
mem[16'h817B] = 8'h58;
mem[16'h817C] = 8'h02;
mem[16'h817D] = 8'h00;
mem[16'h817E] = 8'h3A;
mem[16'h817F] = 8'h70;
mem[16'h8180] = 8'h02;
mem[16'h8181] = 8'h00;
mem[16'h8182] = 8'h3A;
mem[16'h8183] = 8'h70;
mem[16'h8184] = 8'h02;
mem[16'h8185] = 8'h00;
mem[16'h8186] = 8'h3A;
mem[16'h8187] = 8'h70;
mem[16'h8188] = 8'h02;
mem[16'h8189] = 8'h00;
mem[16'h818A] = 8'h6A;
mem[16'h818B] = 8'h58;
mem[16'h818C] = 8'h02;
mem[16'h818D] = 8'h00;
mem[16'h818E] = 8'h00;
mem[16'h818F] = 8'h00;
mem[16'h8190] = 8'h00;
mem[16'h8191] = 8'h00;
mem[16'h8192] = 8'h28;
mem[16'h8193] = 8'h50;
mem[16'h8194] = 8'h00;
mem[16'h8195] = 8'h00;
mem[16'h8196] = 8'h20;
mem[16'h8197] = 8'h10;
mem[16'h8198] = 8'h00;
mem[16'h8199] = 8'h00;
mem[16'h819A] = 8'h40;
mem[16'h819B] = 8'h20;
mem[16'h819C] = 8'h00;
mem[16'h819D] = 8'h00;
mem[16'h819E] = 8'h50;
mem[16'h819F] = 8'h20;
mem[16'h81A0] = 8'h01;
mem[16'h81A1] = 8'h00;
mem[16'h81A2] = 8'h00;
mem[16'h81A3] = 8'h00;
mem[16'h81A4] = 8'h00;
mem[16'h81A5] = 8'h00;
mem[16'h81A6] = 8'h54;
mem[16'h81A7] = 8'h31;
mem[16'h81A8] = 8'h05;
mem[16'h81A9] = 8'h00;
mem[16'h81AA] = 8'h74;
mem[16'h81AB] = 8'h60;
mem[16'h81AC] = 8'h05;
mem[16'h81AD] = 8'h00;
mem[16'h81AE] = 8'h74;
mem[16'h81AF] = 8'h60;
mem[16'h81B0] = 8'h05;
mem[16'h81B1] = 8'h00;
mem[16'h81B2] = 8'h74;
mem[16'h81B3] = 8'h60;
mem[16'h81B4] = 8'h05;
mem[16'h81B5] = 8'h00;
mem[16'h81B6] = 8'h54;
mem[16'h81B7] = 8'h31;
mem[16'h81B8] = 8'h05;
mem[16'h81B9] = 8'h00;
mem[16'h81BA] = 8'h00;
mem[16'h81BB] = 8'h00;
mem[16'h81BC] = 8'h00;
mem[16'h81BD] = 8'h00;
mem[16'h81BE] = 8'h50;
mem[16'h81BF] = 8'h20;
mem[16'h81C0] = 8'h01;
mem[16'h81C1] = 8'h00;
mem[16'h81C2] = 8'h40;
mem[16'h81C3] = 8'h20;
mem[16'h81C4] = 8'h00;
mem[16'h81C5] = 8'h00;
mem[16'h81C6] = 8'h00;
mem[16'h81C7] = 8'h41;
mem[16'h81C8] = 8'h00;
mem[16'h81C9] = 8'h00;
mem[16'h81CA] = 8'h20;
mem[16'h81CB] = 8'h41;
mem[16'h81CC] = 8'h02;
mem[16'h81CD] = 8'h00;
mem[16'h81CE] = 8'h00;
mem[16'h81CF] = 8'h00;
mem[16'h81D0] = 8'h00;
mem[16'h81D1] = 8'h00;
mem[16'h81D2] = 8'h28;
mem[16'h81D3] = 8'h63;
mem[16'h81D4] = 8'h0A;
mem[16'h81D5] = 8'h00;
mem[16'h81D6] = 8'h68;
mem[16'h81D7] = 8'h41;
mem[16'h81D8] = 8'h0B;
mem[16'h81D9] = 8'h00;
mem[16'h81DA] = 8'h68;
mem[16'h81DB] = 8'h41;
mem[16'h81DC] = 8'h0B;
mem[16'h81DD] = 8'h00;
mem[16'h81DE] = 8'h68;
mem[16'h81DF] = 8'h41;
mem[16'h81E0] = 8'h0B;
mem[16'h81E1] = 8'h00;
mem[16'h81E2] = 8'h28;
mem[16'h81E3] = 8'h63;
mem[16'h81E4] = 8'h0A;
mem[16'h81E5] = 8'h00;
mem[16'h81E6] = 8'h00;
mem[16'h81E7] = 8'h00;
mem[16'h81E8] = 8'h00;
mem[16'h81E9] = 8'h00;
mem[16'h81EA] = 8'h20;
mem[16'h81EB] = 8'h41;
mem[16'h81EC] = 8'h02;
mem[16'h81ED] = 8'h00;
mem[16'h81EE] = 8'h00;
mem[16'h81EF] = 8'h41;
mem[16'h81F0] = 8'h00;
mem[16'h81F1] = 8'h00;
mem[16'h81F2] = 8'h00;
mem[16'h81F3] = 8'h02;
mem[16'h81F4] = 8'h01;
mem[16'h81F5] = 8'h00;
mem[16'h81F6] = 8'h40;
mem[16'h81F7] = 8'h02;
mem[16'h81F8] = 8'h05;
mem[16'h81F9] = 8'h00;
mem[16'h81FA] = 8'h00;
mem[16'h81FB] = 8'h00;
mem[16'h81FC] = 8'h00;
mem[16'h81FD] = 8'h00;
mem[16'h81FE] = 8'h50;
mem[16'h81FF] = 8'h46;
mem[16'h8200] = 8'h15;
mem[16'h8201] = 8'h00;
mem[16'h8202] = 8'h50;
mem[16'h8203] = 8'h03;
mem[16'h8204] = 8'h17;
mem[16'h8205] = 8'h00;
mem[16'h8206] = 8'h50;
mem[16'h8207] = 8'h03;
mem[16'h8208] = 8'h17;
mem[16'h8209] = 8'h00;
mem[16'h820A] = 8'h50;
mem[16'h820B] = 8'h03;
mem[16'h820C] = 8'h17;
mem[16'h820D] = 8'h00;
mem[16'h820E] = 8'h50;
mem[16'h820F] = 8'h46;
mem[16'h8210] = 8'h15;
mem[16'h8211] = 8'h00;
mem[16'h8212] = 8'h00;
mem[16'h8213] = 8'h00;
mem[16'h8214] = 8'h00;
mem[16'h8215] = 8'h00;
mem[16'h8216] = 8'h40;
mem[16'h8217] = 8'h02;
mem[16'h8218] = 8'h05;
mem[16'h8219] = 8'h00;
mem[16'h821A] = 8'h00;
mem[16'h821B] = 8'h02;
mem[16'h821C] = 8'h01;
mem[16'h821D] = 8'h00;
mem[16'h821E] = 8'h00;
mem[16'h821F] = 8'h04;
mem[16'h8220] = 8'h02;
mem[16'h8221] = 8'h00;
mem[16'h8222] = 8'h00;
mem[16'h8223] = 8'h05;
mem[16'h8224] = 8'h0A;
mem[16'h8225] = 8'h00;
mem[16'h8226] = 8'h00;
mem[16'h8227] = 8'h00;
mem[16'h8228] = 8'h00;
mem[16'h8229] = 8'h00;
mem[16'h822A] = 8'h20;
mem[16'h822B] = 8'h0D;
mem[16'h822C] = 8'h2B;
mem[16'h822D] = 8'h00;
mem[16'h822E] = 8'h20;
mem[16'h822F] = 8'h07;
mem[16'h8230] = 8'h2E;
mem[16'h8231] = 8'h00;
mem[16'h8232] = 8'h20;
mem[16'h8233] = 8'h07;
mem[16'h8234] = 8'h2E;
mem[16'h8235] = 8'h00;
mem[16'h8236] = 8'h20;
mem[16'h8237] = 8'h07;
mem[16'h8238] = 8'h2E;
mem[16'h8239] = 8'h00;
mem[16'h823A] = 8'h20;
mem[16'h823B] = 8'h0D;
mem[16'h823C] = 8'h2B;
mem[16'h823D] = 8'h00;
mem[16'h823E] = 8'h00;
mem[16'h823F] = 8'h00;
mem[16'h8240] = 8'h00;
mem[16'h8241] = 8'h00;
mem[16'h8242] = 8'h00;
mem[16'h8243] = 8'h05;
mem[16'h8244] = 8'h0A;
mem[16'h8245] = 8'h00;
mem[16'h8246] = 8'h00;
mem[16'h8247] = 8'h04;
mem[16'h8248] = 8'h02;
mem[16'h8249] = 8'h00;
mem[16'h824A] = 8'h00;
mem[16'h824B] = 8'h08;
mem[16'h824C] = 8'h04;
mem[16'h824D] = 8'h00;
mem[16'h824E] = 8'h00;
mem[16'h824F] = 8'h0A;
mem[16'h8250] = 8'h14;
mem[16'h8251] = 8'h00;
mem[16'h8252] = 8'h00;
mem[16'h8253] = 8'h00;
mem[16'h8254] = 8'h00;
mem[16'h8255] = 8'h00;
mem[16'h8256] = 8'h40;
mem[16'h8257] = 8'h1A;
mem[16'h8258] = 8'h56;
mem[16'h8259] = 8'h00;
mem[16'h825A] = 8'h40;
mem[16'h825B] = 8'h0E;
mem[16'h825C] = 8'h5C;
mem[16'h825D] = 8'h00;
mem[16'h825E] = 8'h40;
mem[16'h825F] = 8'h0E;
mem[16'h8260] = 8'h5C;
mem[16'h8261] = 8'h00;
mem[16'h8262] = 8'h40;
mem[16'h8263] = 8'h0E;
mem[16'h8264] = 8'h5C;
mem[16'h8265] = 8'h00;
mem[16'h8266] = 8'h40;
mem[16'h8267] = 8'h1A;
mem[16'h8268] = 8'h56;
mem[16'h8269] = 8'h00;
mem[16'h826A] = 8'h00;
mem[16'h826B] = 8'h00;
mem[16'h826C] = 8'h00;
mem[16'h826D] = 8'h00;
mem[16'h826E] = 8'h00;
mem[16'h826F] = 8'h0A;
mem[16'h8270] = 8'h14;
mem[16'h8271] = 8'h00;
mem[16'h8272] = 8'h00;
mem[16'h8273] = 8'h08;
mem[16'h8274] = 8'h04;
mem[16'h8275] = 8'h00;
mem[16'h8276] = 8'h00;
mem[16'h8277] = 8'h10;
mem[16'h8278] = 8'h08;
mem[16'h8279] = 8'h00;
mem[16'h827A] = 8'h00;
mem[16'h827B] = 8'h14;
mem[16'h827C] = 8'h28;
mem[16'h827D] = 8'h00;
mem[16'h827E] = 8'h00;
mem[16'h827F] = 8'h00;
mem[16'h8280] = 8'h00;
mem[16'h8281] = 8'h00;
mem[16'h8282] = 8'h00;
mem[16'h8283] = 8'h35;
mem[16'h8284] = 8'h2C;
mem[16'h8285] = 8'h01;
mem[16'h8286] = 8'h00;
mem[16'h8287] = 8'h1D;
mem[16'h8288] = 8'h38;
mem[16'h8289] = 8'h01;
mem[16'h828A] = 8'h00;
mem[16'h828B] = 8'h1D;
mem[16'h828C] = 8'h38;
mem[16'h828D] = 8'h01;
mem[16'h828E] = 8'h00;
mem[16'h828F] = 8'h1D;
mem[16'h8290] = 8'h38;
mem[16'h8291] = 8'h01;
mem[16'h8292] = 8'h00;
mem[16'h8293] = 8'h35;
mem[16'h8294] = 8'h2C;
mem[16'h8295] = 8'h01;
mem[16'h8296] = 8'h00;
mem[16'h8297] = 8'h00;
mem[16'h8298] = 8'h00;
mem[16'h8299] = 8'h00;
mem[16'h829A] = 8'h00;
mem[16'h829B] = 8'h14;
mem[16'h829C] = 8'h28;
mem[16'h829D] = 8'h00;
mem[16'h829E] = 8'h00;
mem[16'h829F] = 8'h10;
mem[16'h82A0] = 8'h08;
mem[16'h82A1] = 8'h00;
mem[16'h82A2] = 8'hA0;
mem[16'h82A3] = 8'h00;
mem[16'h82A4] = 8'h8C;
mem[16'h82A5] = 8'h3B;
mem[16'h82A6] = 8'h83;
mem[16'h82A7] = 8'h8C;
mem[16'h82A8] = 8'h3C;
mem[16'h82A9] = 8'h83;
mem[16'h82AA] = 8'h20;
mem[16'h82AB] = 8'hCB;
mem[16'h82AC] = 8'h82;
mem[16'h82AD] = 8'h20;
mem[16'h82AE] = 8'hE4;
mem[16'h82AF] = 8'h82;
mem[16'h82B0] = 8'h20;
mem[16'h82B1] = 8'hF9;
mem[16'h82B2] = 8'h82;
mem[16'h82B3] = 8'hD0;
mem[16'h82B4] = 8'h03;
mem[16'h82B5] = 8'h20;
mem[16'h82B6] = 8'hCB;
mem[16'h82B7] = 8'h82;
mem[16'h82B8] = 8'h20;
mem[16'h82B9] = 8'h1A;
mem[16'h82BA] = 8'h83;
mem[16'h82BB] = 8'hD0;
mem[16'h82BC] = 8'h08;
mem[16'h82BD] = 8'h20;
mem[16'h82BE] = 8'hE4;
mem[16'h82BF] = 8'h82;
mem[16'h82C0] = 8'hA9;
mem[16'h82C1] = 8'hFF;
mem[16'h82C2] = 8'h20;
mem[16'h82C3] = 8'hA8;
mem[16'h82C4] = 8'hFC;
mem[16'h82C5] = 8'h4C;
mem[16'h82C6] = 8'hB0;
mem[16'h82C7] = 8'h82;
mem[16'h82C8] = 8'h68;
mem[16'h82C9] = 8'h68;
mem[16'h82CA] = 8'h60;
mem[16'h82CB] = 8'hAC;
mem[16'h82CC] = 8'h3B;
mem[16'h82CD] = 8'h83;
mem[16'h82CE] = 8'hB1;
mem[16'h82CF] = 8'h79;
mem[16'h82D0] = 8'hC9;
mem[16'h82D1] = 8'hFF;
mem[16'h82D2] = 8'hF0;
mem[16'h82D3] = 8'hF4;
mem[16'h82D4] = 8'h8D;
mem[16'h82D5] = 8'h3D;
mem[16'h82D6] = 8'h83;
mem[16'h82D7] = 8'hC8;
mem[16'h82D8] = 8'hB1;
mem[16'h82D9] = 8'h79;
mem[16'h82DA] = 8'hC8;
mem[16'h82DB] = 8'h4A;
mem[16'h82DC] = 8'h4A;
mem[16'h82DD] = 8'h8D;
mem[16'h82DE] = 8'h3F;
mem[16'h82DF] = 8'h83;
mem[16'h82E0] = 8'h8C;
mem[16'h82E1] = 8'h3B;
mem[16'h82E2] = 8'h83;
mem[16'h82E3] = 8'h60;
mem[16'h82E4] = 8'hAC;
mem[16'h82E5] = 8'h3C;
mem[16'h82E6] = 8'h83;
mem[16'h82E7] = 8'hB1;
mem[16'h82E8] = 8'h7B;
mem[16'h82E9] = 8'h8D;
mem[16'h82EA] = 8'h3E;
mem[16'h82EB] = 8'h83;
mem[16'h82EC] = 8'hC8;
mem[16'h82ED] = 8'hB1;
mem[16'h82EE] = 8'h7B;
mem[16'h82EF] = 8'hC8;
mem[16'h82F0] = 8'h4A;
mem[16'h82F1] = 8'h4A;
mem[16'h82F2] = 8'h8D;
mem[16'h82F3] = 8'h40;
mem[16'h82F4] = 8'h83;
mem[16'h82F5] = 8'h8C;
mem[16'h82F6] = 8'h3C;
mem[16'h82F7] = 8'h83;
mem[16'h82F8] = 8'h60;
mem[16'h82F9] = 8'hAD;
mem[16'h82FA] = 8'h3D;
mem[16'h82FB] = 8'h83;
mem[16'h82FC] = 8'hD0;
mem[16'h82FD] = 8'h09;
mem[16'h82FE] = 8'hA9;
mem[16'h82FF] = 8'h96;
mem[16'h8300] = 8'h20;
mem[16'h8301] = 8'hA8;
mem[16'h8302] = 8'hFC;
mem[16'h8303] = 8'hCE;
mem[16'h8304] = 8'h3F;
mem[16'h8305] = 8'h83;
mem[16'h8306] = 8'h60;
mem[16'h8307] = 8'h85;
mem[16'h8308] = 8'h50;
mem[16'h8309] = 8'hA9;
mem[16'h830A] = 8'h0A;
mem[16'h830B] = 8'h85;
mem[16'h830C] = 8'h52;
mem[16'h830D] = 8'h85;
mem[16'h830E] = 8'h53;
mem[16'h830F] = 8'hA9;
mem[16'h8310] = 8'h00;
mem[16'h8311] = 8'h85;
mem[16'h8312] = 8'h55;
mem[16'h8313] = 8'h20;
mem[16'h8314] = 8'h00;
mem[16'h8315] = 8'h65;
mem[16'h8316] = 8'hCE;
mem[16'h8317] = 8'h3F;
mem[16'h8318] = 8'h83;
mem[16'h8319] = 8'h60;
mem[16'h831A] = 8'hAD;
mem[16'h831B] = 8'h3E;
mem[16'h831C] = 8'h83;
mem[16'h831D] = 8'hD0;
mem[16'h831E] = 8'h09;
mem[16'h831F] = 8'hA9;
mem[16'h8320] = 8'hFF;
mem[16'h8321] = 8'h20;
mem[16'h8322] = 8'hA8;
mem[16'h8323] = 8'hFC;
mem[16'h8324] = 8'hCE;
mem[16'h8325] = 8'h40;
mem[16'h8326] = 8'h83;
mem[16'h8327] = 8'h60;
mem[16'h8328] = 8'h85;
mem[16'h8329] = 8'h50;
mem[16'h832A] = 8'hA9;
mem[16'h832B] = 8'h06;
mem[16'h832C] = 8'h85;
mem[16'h832D] = 8'h52;
mem[16'h832E] = 8'h85;
mem[16'h832F] = 8'h53;
mem[16'h8330] = 8'hA9;
mem[16'h8331] = 8'h00;
mem[16'h8332] = 8'h85;
mem[16'h8333] = 8'h55;
mem[16'h8334] = 8'h20;
mem[16'h8335] = 8'h00;
mem[16'h8336] = 8'h65;
mem[16'h8337] = 8'hCE;
mem[16'h8338] = 8'h40;
mem[16'h8339] = 8'h83;
mem[16'h833A] = 8'h60;
mem[16'h833B] = 8'h06;
mem[16'h833C] = 8'h04;
mem[16'h833D] = 8'h18;
mem[16'h833E] = 8'h26;
mem[16'h833F] = 8'h01;
mem[16'h8340] = 8'h01;
mem[16'h8341] = 8'h13;
mem[16'h8342] = 8'h04;
mem[16'h8343] = 8'h18;
mem[16'h8344] = 8'h04;
mem[16'h8345] = 8'h18;
mem[16'h8346] = 8'h04;
mem[16'h8347] = 8'h18;
mem[16'h8348] = 8'h04;
mem[16'h8349] = 8'h13;
mem[16'h834A] = 8'h04;
mem[16'h834B] = 8'h18;
mem[16'h834C] = 8'h04;
mem[16'h834D] = 8'h18;
mem[16'h834E] = 8'h04;
mem[16'h834F] = 8'h18;
mem[16'h8350] = 8'h04;
mem[16'h8351] = 8'h12;
mem[16'h8352] = 8'h04;
mem[16'h8353] = 8'h12;
mem[16'h8354] = 8'h04;
mem[16'h8355] = 8'h13;
mem[16'h8356] = 8'h04;
mem[16'h8357] = 8'h13;
mem[16'h8358] = 8'h04;
mem[16'h8359] = 8'h15;
mem[16'h835A] = 8'h04;
mem[16'h835B] = 8'h15;
mem[16'h835C] = 8'h04;
mem[16'h835D] = 8'h00;
mem[16'h835E] = 8'h04;
mem[16'h835F] = 8'h00;
mem[16'h8360] = 8'h04;
mem[16'h8361] = 8'h12;
mem[16'h8362] = 8'h04;
mem[16'h8363] = 8'h12;
mem[16'h8364] = 8'h04;
mem[16'h8365] = 8'h13;
mem[16'h8366] = 8'h04;
mem[16'h8367] = 8'h13;
mem[16'h8368] = 8'h04;
mem[16'h8369] = 8'h15;
mem[16'h836A] = 8'h04;
mem[16'h836B] = 8'h15;
mem[16'h836C] = 8'h04;
mem[16'h836D] = 8'h0E;
mem[16'h836E] = 8'h04;
mem[16'h836F] = 8'h0E;
mem[16'h8370] = 8'h04;
mem[16'h8371] = 8'h10;
mem[16'h8372] = 8'h04;
mem[16'h8373] = 8'h12;
mem[16'h8374] = 8'h04;
mem[16'h8375] = 8'h13;
mem[16'h8376] = 8'h04;
mem[16'h8377] = 8'h15;
mem[16'h8378] = 8'h04;
mem[16'h8379] = 8'h18;
mem[16'h837A] = 8'h08;
mem[16'h837B] = 8'h00;
mem[16'h837C] = 8'h08;
mem[16'h837D] = 8'hFF;
mem[16'h837E] = 8'h30;
mem[16'h837F] = 8'h04;
mem[16'h8380] = 8'h26;
mem[16'h8381] = 8'h04;
mem[16'h8382] = 8'h41;
mem[16'h8383] = 8'h04;
mem[16'h8384] = 8'h26;
mem[16'h8385] = 8'h04;
mem[16'h8386] = 8'h30;
mem[16'h8387] = 8'h04;
mem[16'h8388] = 8'h26;
mem[16'h8389] = 8'h04;
mem[16'h838A] = 8'h41;
mem[16'h838B] = 8'h04;
mem[16'h838C] = 8'h26;
mem[16'h838D] = 8'h04;
mem[16'h838E] = 8'h2B;
mem[16'h838F] = 8'h04;
mem[16'h8390] = 8'h24;
mem[16'h8391] = 8'h04;
mem[16'h8392] = 8'h39;
mem[16'h8393] = 8'h04;
mem[16'h8394] = 8'h24;
mem[16'h8395] = 8'h04;
mem[16'h8396] = 8'h2B;
mem[16'h8397] = 8'h04;
mem[16'h8398] = 8'h24;
mem[16'h8399] = 8'h04;
mem[16'h839A] = 8'h39;
mem[16'h839B] = 8'h04;
mem[16'h839C] = 8'h00;
mem[16'h839D] = 8'h04;
mem[16'h839E] = 8'h2B;
mem[16'h839F] = 8'h04;
mem[16'h83A0] = 8'h24;
mem[16'h83A1] = 8'h04;
mem[16'h83A2] = 8'h39;
mem[16'h83A3] = 8'h04;
mem[16'h83A4] = 8'h24;
mem[16'h83A5] = 8'h04;
mem[16'h83A6] = 8'h2B;
mem[16'h83A7] = 8'h04;
mem[16'h83A8] = 8'h24;
mem[16'h83A9] = 8'h04;
mem[16'h83AA] = 8'h39;
mem[16'h83AB] = 8'h04;
mem[16'h83AC] = 8'h24;
mem[16'h83AD] = 8'h04;
mem[16'h83AE] = 8'h2B;
mem[16'h83AF] = 8'h04;
mem[16'h83B0] = 8'h20;
mem[16'h83B1] = 8'h04;
mem[16'h83B2] = 8'h33;
mem[16'h83B3] = 8'h04;
mem[16'h83B4] = 8'h20;
mem[16'h83B5] = 8'h04;
mem[16'h83B6] = 8'h30;
mem[16'h83B7] = 8'h08;
mem[16'h83B8] = 8'h00;
mem[16'h83B9] = 8'h08;
mem[16'h83BA] = 8'h18;
mem[16'h83BB] = 8'h04;
mem[16'h83BC] = 8'h15;
mem[16'h83BD] = 8'h04;
mem[16'h83BE] = 8'h13;
mem[16'h83BF] = 8'h04;
mem[16'h83C0] = 8'h12;
mem[16'h83C1] = 8'h04;
mem[16'h83C2] = 8'h10;
mem[16'h83C3] = 8'h04;
mem[16'h83C4] = 8'h10;
mem[16'h83C5] = 8'h04;
mem[16'h83C6] = 8'h13;
mem[16'h83C7] = 8'h04;
mem[16'h83C8] = 8'h13;
mem[16'h83C9] = 8'h04;
mem[16'h83CA] = 8'h18;
mem[16'h83CB] = 8'h04;
mem[16'h83CC] = 8'h15;
mem[16'h83CD] = 8'h04;
mem[16'h83CE] = 8'h13;
mem[16'h83CF] = 8'h04;
mem[16'h83D0] = 8'h15;
mem[16'h83D1] = 8'h04;
mem[16'h83D2] = 8'h18;
mem[16'h83D3] = 8'h04;
mem[16'h83D4] = 8'h18;
mem[16'h83D5] = 8'h04;
mem[16'h83D6] = 8'h18;
mem[16'h83D7] = 8'h04;
mem[16'h83D8] = 8'h18;
mem[16'h83D9] = 8'h04;
mem[16'h83DA] = 8'h18;
mem[16'h83DB] = 8'h04;
mem[16'h83DC] = 8'h15;
mem[16'h83DD] = 8'h04;
mem[16'h83DE] = 8'h13;
mem[16'h83DF] = 8'h04;
mem[16'h83E0] = 8'h12;
mem[16'h83E1] = 8'h04;
mem[16'h83E2] = 8'h10;
mem[16'h83E3] = 8'h04;
mem[16'h83E4] = 8'h10;
mem[16'h83E5] = 8'h04;
mem[16'h83E6] = 8'h13;
mem[16'h83E7] = 8'h04;
mem[16'h83E8] = 8'h13;
mem[16'h83E9] = 8'h04;
mem[16'h83EA] = 8'h10;
mem[16'h83EB] = 8'h04;
mem[16'h83EC] = 8'h12;
mem[16'h83ED] = 8'h04;
mem[16'h83EE] = 8'h13;
mem[16'h83EF] = 8'h04;
mem[16'h83F0] = 8'h15;
mem[16'h83F1] = 8'h04;
mem[16'h83F2] = 8'h18;
mem[16'h83F3] = 8'h04;
mem[16'h83F4] = 8'h18;
mem[16'h83F5] = 8'h04;
mem[16'h83F6] = 8'h00;
mem[16'h83F7] = 8'h04;
mem[16'h83F8] = 8'h00;
mem[16'h83F9] = 8'h04;
mem[16'h83FA] = 8'hFF;
mem[16'h83FB] = 8'h30;
mem[16'h83FC] = 8'h04;
mem[16'h83FD] = 8'h26;
mem[16'h83FE] = 8'h04;
mem[16'h83FF] = 8'h30;
mem[16'h8400] = 8'h04;
mem[16'h8401] = 8'h26;
mem[16'h8402] = 8'h04;
mem[16'h8403] = 8'h30;
mem[16'h8404] = 8'h04;
mem[16'h8405] = 8'h26;
mem[16'h8406] = 8'h04;
mem[16'h8407] = 8'h30;
mem[16'h8408] = 8'h04;
mem[16'h8409] = 8'h26;
mem[16'h840A] = 8'h04;
mem[16'h840B] = 8'h30;
mem[16'h840C] = 8'h04;
mem[16'h840D] = 8'h26;
mem[16'h840E] = 8'h04;
mem[16'h840F] = 8'h30;
mem[16'h8410] = 8'h04;
mem[16'h8411] = 8'h26;
mem[16'h8412] = 8'h04;
mem[16'h8413] = 8'h30;
mem[16'h8414] = 8'h04;
mem[16'h8415] = 8'h26;
mem[16'h8416] = 8'h04;
mem[16'h8417] = 8'h30;
mem[16'h8418] = 8'h04;
mem[16'h8419] = 8'h26;
mem[16'h841A] = 8'h04;
mem[16'h841B] = 8'h30;
mem[16'h841C] = 8'h04;
mem[16'h841D] = 8'h26;
mem[16'h841E] = 8'h04;
mem[16'h841F] = 8'h30;
mem[16'h8420] = 8'h04;
mem[16'h8421] = 8'h26;
mem[16'h8422] = 8'h04;
mem[16'h8423] = 8'h30;
mem[16'h8424] = 8'h04;
mem[16'h8425] = 8'h26;
mem[16'h8426] = 8'h04;
mem[16'h8427] = 8'h30;
mem[16'h8428] = 8'h04;
mem[16'h8429] = 8'h26;
mem[16'h842A] = 8'h04;
mem[16'h842B] = 8'h2B;
mem[16'h842C] = 8'h04;
mem[16'h842D] = 8'h20;
mem[16'h842E] = 8'h04;
mem[16'h842F] = 8'h2B;
mem[16'h8430] = 8'h04;
mem[16'h8431] = 8'h20;
mem[16'h8432] = 8'h04;
mem[16'h8433] = 8'h30;
mem[16'h8434] = 8'h04;
mem[16'h8435] = 8'h30;
mem[16'h8436] = 8'h04;
mem[16'h8437] = 8'h00;
mem[16'h8438] = 8'h04;
mem[16'h8439] = 8'h00;
mem[16'h843A] = 8'h04;
mem[16'h843B] = 8'h00;
mem[16'h843C] = 8'h00;
mem[16'h843D] = 8'h00;
mem[16'h843E] = 8'h00;
mem[16'h843F] = 8'h00;
mem[16'h8440] = 8'h00;
mem[16'h8441] = 8'h00;
mem[16'h8442] = 8'h00;
mem[16'h8443] = 8'h20;
mem[16'h8444] = 8'h10;
mem[16'h8445] = 8'h00;
mem[16'h8446] = 8'h00;
mem[16'h8447] = 8'h00;
mem[16'h8448] = 8'h00;
mem[16'h8449] = 8'h00;
mem[16'h844A] = 8'h00;
mem[16'h844B] = 8'h68;
mem[16'h844C] = 8'h5D;
mem[16'h844D] = 8'h00;
mem[16'h844E] = 8'h00;
mem[16'h844F] = 8'h48;
mem[16'h8450] = 8'h48;
mem[16'h8451] = 8'h00;
mem[16'h8452] = 8'h00;
mem[16'h8453] = 8'h68;
mem[16'h8454] = 8'h5D;
mem[16'h8455] = 8'h00;
mem[16'h8456] = 8'h00;
mem[16'h8457] = 8'h00;
mem[16'h8458] = 8'h00;
mem[16'h8459] = 8'h00;
mem[16'h845A] = 8'h00;
mem[16'h845B] = 8'h20;
mem[16'h845C] = 8'h10;
mem[16'h845D] = 8'h00;
mem[16'h845E] = 8'h00;
mem[16'h845F] = 8'h00;
mem[16'h8460] = 8'h00;
mem[16'h8461] = 8'h00;
mem[16'h8462] = 8'h00;
mem[16'h8463] = 8'h00;
mem[16'h8464] = 8'h00;
mem[16'h8465] = 8'h00;
mem[16'h8466] = 8'h00;
mem[16'h8467] = 8'h40;
mem[16'h8468] = 8'h20;
mem[16'h8469] = 8'h00;
mem[16'h846A] = 8'h00;
mem[16'h846B] = 8'h00;
mem[16'h846C] = 8'h00;
mem[16'h846D] = 8'h00;
mem[16'h846E] = 8'h00;
mem[16'h846F] = 8'h50;
mem[16'h8470] = 8'h3B;
mem[16'h8471] = 8'h01;
mem[16'h8472] = 8'h00;
mem[16'h8473] = 8'h10;
mem[16'h8474] = 8'h11;
mem[16'h8475] = 8'h01;
mem[16'h8476] = 8'h00;
mem[16'h8477] = 8'h50;
mem[16'h8478] = 8'h3B;
mem[16'h8479] = 8'h01;
mem[16'h847A] = 8'h00;
mem[16'h847B] = 8'h00;
mem[16'h847C] = 8'h00;
mem[16'h847D] = 8'h00;
mem[16'h847E] = 8'h00;
mem[16'h847F] = 8'h40;
mem[16'h8480] = 8'h20;
mem[16'h8481] = 8'h00;
mem[16'h8482] = 8'h00;
mem[16'h8483] = 8'h00;
mem[16'h8484] = 8'h00;
mem[16'h8485] = 8'h00;
mem[16'h8486] = 8'h00;
mem[16'h8487] = 8'h00;
mem[16'h8488] = 8'h00;
mem[16'h8489] = 8'h00;
mem[16'h848A] = 8'h00;
mem[16'h848B] = 8'h00;
mem[16'h848C] = 8'h41;
mem[16'h848D] = 8'h00;
mem[16'h848E] = 8'h00;
mem[16'h848F] = 8'h00;
mem[16'h8490] = 8'h00;
mem[16'h8491] = 8'h00;
mem[16'h8492] = 8'h00;
mem[16'h8493] = 8'h20;
mem[16'h8494] = 8'h77;
mem[16'h8495] = 8'h02;
mem[16'h8496] = 8'h00;
mem[16'h8497] = 8'h20;
mem[16'h8498] = 8'h22;
mem[16'h8499] = 8'h02;
mem[16'h849A] = 8'h00;
mem[16'h849B] = 8'h20;
mem[16'h849C] = 8'h77;
mem[16'h849D] = 8'h02;
mem[16'h849E] = 8'h00;
mem[16'h849F] = 8'h00;
mem[16'h84A0] = 8'h00;
mem[16'h84A1] = 8'h00;
mem[16'h84A2] = 8'h00;
mem[16'h84A3] = 8'h00;
mem[16'h84A4] = 8'h41;
mem[16'h84A5] = 8'h00;
mem[16'h84A6] = 8'h00;
mem[16'h84A7] = 8'h00;
mem[16'h84A8] = 8'h00;
mem[16'h84A9] = 8'h00;
mem[16'h84AA] = 8'h00;
mem[16'h84AB] = 8'h00;
mem[16'h84AC] = 8'h00;
mem[16'h84AD] = 8'h00;
mem[16'h84AE] = 8'h00;
mem[16'h84AF] = 8'h00;
mem[16'h84B0] = 8'h02;
mem[16'h84B1] = 8'h01;
mem[16'h84B2] = 8'h00;
mem[16'h84B3] = 8'h00;
mem[16'h84B4] = 8'h00;
mem[16'h84B5] = 8'h00;
mem[16'h84B6] = 8'h00;
mem[16'h84B7] = 8'h40;
mem[16'h84B8] = 8'h6E;
mem[16'h84B9] = 8'h05;
mem[16'h84BA] = 8'h00;
mem[16'h84BB] = 8'h40;
mem[16'h84BC] = 8'h44;
mem[16'h84BD] = 8'h04;
mem[16'h84BE] = 8'h00;
mem[16'h84BF] = 8'h40;
mem[16'h84C0] = 8'h6E;
mem[16'h84C1] = 8'h05;
mem[16'h84C2] = 8'h00;
mem[16'h84C3] = 8'h00;
mem[16'h84C4] = 8'h00;
mem[16'h84C5] = 8'h00;
mem[16'h84C6] = 8'h00;
mem[16'h84C7] = 8'h00;
mem[16'h84C8] = 8'h02;
mem[16'h84C9] = 8'h01;
mem[16'h84CA] = 8'h00;
mem[16'h84CB] = 8'h00;
mem[16'h84CC] = 8'h00;
mem[16'h84CD] = 8'h00;
mem[16'h84CE] = 8'h00;
mem[16'h84CF] = 8'h00;
mem[16'h84D0] = 8'h00;
mem[16'h84D1] = 8'h00;
mem[16'h84D2] = 8'h00;
mem[16'h84D3] = 8'h00;
mem[16'h84D4] = 8'h04;
mem[16'h84D5] = 8'h02;
mem[16'h84D6] = 8'h00;
mem[16'h84D7] = 8'h00;
mem[16'h84D8] = 8'h00;
mem[16'h84D9] = 8'h00;
mem[16'h84DA] = 8'h00;
mem[16'h84DB] = 8'h00;
mem[16'h84DC] = 8'h5D;
mem[16'h84DD] = 8'h0B;
mem[16'h84DE] = 8'h00;
mem[16'h84DF] = 8'h00;
mem[16'h84E0] = 8'h09;
mem[16'h84E1] = 8'h09;
mem[16'h84E2] = 8'h00;
mem[16'h84E3] = 8'h00;
mem[16'h84E4] = 8'h5D;
mem[16'h84E5] = 8'h0B;
mem[16'h84E6] = 8'h00;
mem[16'h84E7] = 8'h00;
mem[16'h84E8] = 8'h00;
mem[16'h84E9] = 8'h00;
mem[16'h84EA] = 8'h00;
mem[16'h84EB] = 8'h00;
mem[16'h84EC] = 8'h04;
mem[16'h84ED] = 8'h02;
mem[16'h84EE] = 8'h00;
mem[16'h84EF] = 8'h00;
mem[16'h84F0] = 8'h00;
mem[16'h84F1] = 8'h00;
mem[16'h84F2] = 8'h00;
mem[16'h84F3] = 8'h00;
mem[16'h84F4] = 8'h00;
mem[16'h84F5] = 8'h00;
mem[16'h84F6] = 8'h00;
mem[16'h84F7] = 8'h00;
mem[16'h84F8] = 8'h08;
mem[16'h84F9] = 8'h04;
mem[16'h84FA] = 8'h00;
mem[16'h84FB] = 8'h00;
mem[16'h84FC] = 8'h00;
mem[16'h84FD] = 8'h00;
mem[16'h84FE] = 8'h00;
mem[16'h84FF] = 8'h00;
mem[16'h8500] = 8'h3A;
mem[16'h8501] = 8'h17;
mem[16'h8502] = 8'h00;
mem[16'h8503] = 8'h00;
mem[16'h8504] = 8'h12;
mem[16'h8505] = 8'h12;
mem[16'h8506] = 8'h00;
mem[16'h8507] = 8'h00;
mem[16'h8508] = 8'h3A;
mem[16'h8509] = 8'h17;
mem[16'h850A] = 8'h00;
mem[16'h850B] = 8'h00;
mem[16'h850C] = 8'h00;
mem[16'h850D] = 8'h00;
mem[16'h850E] = 8'h00;
mem[16'h850F] = 8'h00;
mem[16'h8510] = 8'h08;
mem[16'h8511] = 8'h04;
mem[16'h8512] = 8'h00;
mem[16'h8513] = 8'h00;
mem[16'h8514] = 8'h00;
mem[16'h8515] = 8'h00;
mem[16'h8516] = 8'h00;
mem[16'h8517] = 8'h00;
mem[16'h8518] = 8'h00;
mem[16'h8519] = 8'h00;
mem[16'h851A] = 8'h00;
mem[16'h851B] = 8'h00;
mem[16'h851C] = 8'h10;
mem[16'h851D] = 8'h08;
mem[16'h851E] = 8'h00;
mem[16'h851F] = 8'h00;
mem[16'h8520] = 8'h00;
mem[16'h8521] = 8'h00;
mem[16'h8522] = 8'h00;
mem[16'h8523] = 8'h00;
mem[16'h8524] = 8'h74;
mem[16'h8525] = 8'h2E;
mem[16'h8526] = 8'h00;
mem[16'h8527] = 8'h00;
mem[16'h8528] = 8'h24;
mem[16'h8529] = 8'h24;
mem[16'h852A] = 8'h00;
mem[16'h852B] = 8'h00;
mem[16'h852C] = 8'h74;
mem[16'h852D] = 8'h2E;
mem[16'h852E] = 8'h00;
mem[16'h852F] = 8'h00;
mem[16'h8530] = 8'h00;
mem[16'h8531] = 8'h00;
mem[16'h8532] = 8'h00;
mem[16'h8533] = 8'h00;
mem[16'h8534] = 8'h10;
mem[16'h8535] = 8'h08;
mem[16'h8536] = 8'h00;
mem[16'h8537] = 8'hAD;
mem[16'h8538] = 8'hAF;
mem[16'h8539] = 8'h85;
mem[16'h853A] = 8'h85;
mem[16'h853B] = 8'h56;
mem[16'h853C] = 8'hA9;
mem[16'h853D] = 8'h51;
mem[16'h853E] = 8'hA0;
mem[16'h853F] = 8'h85;
mem[16'h8540] = 8'h20;
mem[16'h8541] = 8'h2B;
mem[16'h8542] = 8'h8C;
mem[16'h8543] = 8'hA9;
mem[16'h8544] = 8'h12;
mem[16'h8545] = 8'h8D;
mem[16'h8546] = 8'h24;
mem[16'h8547] = 8'h8C;
mem[16'h8548] = 8'hAD;
mem[16'h8549] = 8'hAE;
mem[16'h854A] = 8'h85;
mem[16'h854B] = 8'h85;
mem[16'h854C] = 8'h57;
mem[16'h854D] = 8'h20;
mem[16'h854E] = 8'hA8;
mem[16'h854F] = 8'h8B;
mem[16'h8550] = 8'h60;
mem[16'h8551] = 8'h00;
mem[16'h8552] = 8'h30;
mem[16'h8553] = 8'h1B;
mem[16'h8554] = 8'h0C;
mem[16'h8555] = 8'h27;
mem[16'h8556] = 8'h3F;
mem[16'h8557] = 8'h2C;
mem[16'h8558] = 8'h35;
mem[16'h8559] = 8'h2C;
mem[16'h855A] = 8'h35;
mem[16'h855B] = 8'h2C;
mem[16'h855C] = 8'h35;
mem[16'h855D] = 8'h27;
mem[16'h855E] = 8'h3F;
mem[16'h855F] = 8'h1B;
mem[16'h8560] = 8'h0C;
mem[16'h8561] = 8'h00;
mem[16'h8562] = 8'h30;
mem[16'h8563] = 8'hAD;
mem[16'h8564] = 8'hB0;
mem[16'h8565] = 8'h85;
mem[16'h8566] = 8'hD0;
mem[16'h8567] = 8'h45;
mem[16'h8568] = 8'hAD;
mem[16'h8569] = 8'hB2;
mem[16'h856A] = 8'h85;
mem[16'h856B] = 8'hD0;
mem[16'h856C] = 8'h40;
mem[16'h856D] = 8'hAD;
mem[16'h856E] = 8'h13;
mem[16'h856F] = 8'h87;
mem[16'h8570] = 8'h29;
mem[16'h8571] = 8'h01;
mem[16'h8572] = 8'hAA;
mem[16'h8573] = 8'hBD;
mem[16'h8574] = 8'h1F;
mem[16'h8575] = 8'h53;
mem[16'h8576] = 8'hC9;
mem[16'h8577] = 8'hFA;
mem[16'h8578] = 8'hB0;
mem[16'h8579] = 8'h33;
mem[16'h857A] = 8'hC9;
mem[16'h857B] = 8'h20;
mem[16'h857C] = 8'h90;
mem[16'h857D] = 8'h2F;
mem[16'h857E] = 8'h38;
mem[16'h857F] = 8'hE9;
mem[16'h8580] = 8'h1E;
mem[16'h8581] = 8'h90;
mem[16'h8582] = 8'h2A;
mem[16'h8583] = 8'h8D;
mem[16'h8584] = 8'hAE;
mem[16'h8585] = 8'h85;
mem[16'h8586] = 8'hAD;
mem[16'h8587] = 8'hD0;
mem[16'h8588] = 8'h4D;
mem[16'h8589] = 8'hC9;
mem[16'h858A] = 8'h3F;
mem[16'h858B] = 8'hD0;
mem[16'h858C] = 8'h0E;
mem[16'h858D] = 8'hAD;
mem[16'h858E] = 8'hCF;
mem[16'h858F] = 8'h4D;
mem[16'h8590] = 8'h38;
mem[16'h8591] = 8'hED;
mem[16'h8592] = 8'hAE;
mem[16'h8593] = 8'h85;
mem[16'h8594] = 8'h20;
mem[16'h8595] = 8'h62;
mem[16'h8596] = 8'h65;
mem[16'h8597] = 8'hC9;
mem[16'h8598] = 8'h0E;
mem[16'h8599] = 8'h90;
mem[16'h859A] = 8'h12;
mem[16'h859B] = 8'hA9;
mem[16'h859C] = 8'h41;
mem[16'h859D] = 8'h8D;
mem[16'h859E] = 8'hAF;
mem[16'h859F] = 8'h85;
mem[16'h85A0] = 8'h20;
mem[16'h85A1] = 8'h37;
mem[16'h85A2] = 8'h85;
mem[16'h85A3] = 8'hA9;
mem[16'h85A4] = 8'h01;
mem[16'h85A5] = 8'h8D;
mem[16'h85A6] = 8'hB2;
mem[16'h85A7] = 8'h85;
mem[16'h85A8] = 8'hA9;
mem[16'h85A9] = 8'h00;
mem[16'h85AA] = 8'h8D;
mem[16'h85AB] = 8'hB3;
mem[16'h85AC] = 8'h85;
mem[16'h85AD] = 8'h60;
mem[16'h85AE] = 8'h20;
mem[16'h85AF] = 8'hC4;
mem[16'h85B0] = 8'h46;
mem[16'h85B1] = 8'h46;
mem[16'h85B2] = 8'h00;
mem[16'h85B3] = 8'h00;
mem[16'h85B4] = 8'hAD;
mem[16'h85B5] = 8'hB2;
mem[16'h85B6] = 8'h85;
mem[16'h85B7] = 8'hF0;
mem[16'h85B8] = 8'h1D;
mem[16'h85B9] = 8'h20;
mem[16'h85BA] = 8'hD7;
mem[16'h85BB] = 8'h85;
mem[16'h85BC] = 8'hAD;
mem[16'h85BD] = 8'hAE;
mem[16'h85BE] = 8'h85;
mem[16'h85BF] = 8'h18;
mem[16'h85C0] = 8'h69;
mem[16'h85C1] = 8'h02;
mem[16'h85C2] = 8'h8D;
mem[16'h85C3] = 8'hAE;
mem[16'h85C4] = 8'h85;
mem[16'h85C5] = 8'hC9;
mem[16'h85C6] = 8'hEA;
mem[16'h85C7] = 8'h90;
mem[16'h85C8] = 8'h0D;
mem[16'h85C9] = 8'h20;
mem[16'h85CA] = 8'h37;
mem[16'h85CB] = 8'h85;
mem[16'h85CC] = 8'hA9;
mem[16'h85CD] = 8'hFF;
mem[16'h85CE] = 8'h8D;
mem[16'h85CF] = 8'hB0;
mem[16'h85D0] = 8'h85;
mem[16'h85D1] = 8'hA9;
mem[16'h85D2] = 8'h00;
mem[16'h85D3] = 8'h8D;
mem[16'h85D4] = 8'hB2;
mem[16'h85D5] = 8'h85;
mem[16'h85D6] = 8'h60;
mem[16'h85D7] = 8'hAD;
mem[16'h85D8] = 8'hAF;
mem[16'h85D9] = 8'h85;
mem[16'h85DA] = 8'h85;
mem[16'h85DB] = 8'h56;
mem[16'h85DC] = 8'hAC;
mem[16'h85DD] = 8'hAE;
mem[16'h85DE] = 8'h85;
mem[16'h85DF] = 8'h84;
mem[16'h85E0] = 8'h57;
mem[16'h85E1] = 8'hB9;
mem[16'h85E2] = 8'h3E;
mem[16'h85E3] = 8'h8C;
mem[16'h85E4] = 8'hAA;
mem[16'h85E5] = 8'hBD;
mem[16'h85E6] = 8'h94;
mem[16'h85E7] = 8'h8E;
mem[16'h85E8] = 8'hAA;
mem[16'h85E9] = 8'hBD;
mem[16'h85EA] = 8'h31;
mem[16'h85EB] = 8'h86;
mem[16'h85EC] = 8'hBC;
mem[16'h85ED] = 8'h38;
mem[16'h85EE] = 8'h86;
mem[16'h85EF] = 8'h20;
mem[16'h85F0] = 8'h3B;
mem[16'h85F1] = 8'h8B;
mem[16'h85F2] = 8'hA9;
mem[16'h85F3] = 8'h1B;
mem[16'h85F4] = 8'h8D;
mem[16'h85F5] = 8'h34;
mem[16'h85F6] = 8'h8B;
mem[16'h85F7] = 8'h20;
mem[16'h85F8] = 8'hF0;
mem[16'h85F9] = 8'h8A;
mem[16'h85FA] = 8'h60;
mem[16'h85FB] = 8'hAD;
mem[16'h85FC] = 8'hB2;
mem[16'h85FD] = 8'h85;
mem[16'h85FE] = 8'hF0;
mem[16'h85FF] = 8'h30;
mem[16'h8600] = 8'hAD;
mem[16'h8601] = 8'hD0;
mem[16'h8602] = 8'h4D;
mem[16'h8603] = 8'hC9;
mem[16'h8604] = 8'h3F;
mem[16'h8605] = 8'hD0;
mem[16'h8606] = 8'h29;
mem[16'h8607] = 8'hAD;
mem[16'h8608] = 8'hCF;
mem[16'h8609] = 8'h4D;
mem[16'h860A] = 8'h38;
mem[16'h860B] = 8'hED;
mem[16'h860C] = 8'hAE;
mem[16'h860D] = 8'h85;
mem[16'h860E] = 8'h20;
mem[16'h860F] = 8'h62;
mem[16'h8610] = 8'h65;
mem[16'h8611] = 8'hC9;
mem[16'h8612] = 8'h0C;
mem[16'h8613] = 8'hB0;
mem[16'h8614] = 8'h1B;
mem[16'h8615] = 8'hA9;
mem[16'h8616] = 8'h01;
mem[16'h8617] = 8'h8D;
mem[16'h8618] = 8'hB3;
mem[16'h8619] = 8'h85;
mem[16'h861A] = 8'h20;
mem[16'h861B] = 8'hAE;
mem[16'h861C] = 8'h4C;
mem[16'h861D] = 8'h20;
mem[16'h861E] = 8'h37;
mem[16'h861F] = 8'h85;
mem[16'h8620] = 8'h20;
mem[16'h8621] = 8'hAE;
mem[16'h8622] = 8'h4C;
mem[16'h8623] = 8'hA9;
mem[16'h8624] = 8'hFF;
mem[16'h8625] = 8'h8D;
mem[16'h8626] = 8'hB0;
mem[16'h8627] = 8'h85;
mem[16'h8628] = 8'hA9;
mem[16'h8629] = 8'h00;
mem[16'h862A] = 8'h8D;
mem[16'h862B] = 8'hB2;
mem[16'h862C] = 8'h85;
mem[16'h862D] = 8'h20;
mem[16'h862E] = 8'h0E;
mem[16'h862F] = 8'h73;
mem[16'h8630] = 8'h60;
mem[16'h8631] = 8'h3F;
mem[16'h8632] = 8'h5A;
mem[16'h8633] = 8'h75;
mem[16'h8634] = 8'h90;
mem[16'h8635] = 8'hAB;
mem[16'h8636] = 8'hC6;
mem[16'h8637] = 8'hE1;
mem[16'h8638] = 8'h86;
mem[16'h8639] = 8'h86;
mem[16'h863A] = 8'h86;
mem[16'h863B] = 8'h86;
mem[16'h863C] = 8'h86;
mem[16'h863D] = 8'h86;
mem[16'h863E] = 8'h86;
mem[16'h863F] = 8'h00;
mem[16'h8640] = 8'h70;
mem[16'h8641] = 8'h01;
mem[16'h8642] = 8'h77;
mem[16'h8643] = 8'h3C;
mem[16'h8644] = 8'h00;
mem[16'h8645] = 8'h3B;
mem[16'h8646] = 8'h42;
mem[16'h8647] = 8'h01;
mem[16'h8648] = 8'h1C;
mem[16'h8649] = 8'h60;
mem[16'h864A] = 8'h01;
mem[16'h864B] = 8'h1C;
mem[16'h864C] = 8'h60;
mem[16'h864D] = 8'h01;
mem[16'h864E] = 8'h1C;
mem[16'h864F] = 8'h60;
mem[16'h8650] = 8'h01;
mem[16'h8651] = 8'h3B;
mem[16'h8652] = 8'h42;
mem[16'h8653] = 8'h01;
mem[16'h8654] = 8'h77;
mem[16'h8655] = 8'h3C;
mem[16'h8656] = 8'h00;
mem[16'h8657] = 8'h00;
mem[16'h8658] = 8'h70;
mem[16'h8659] = 8'h01;
mem[16'h865A] = 8'h00;
mem[16'h865B] = 8'h60;
mem[16'h865C] = 8'h03;
mem[16'h865D] = 8'h6E;
mem[16'h865E] = 8'h79;
mem[16'h865F] = 8'h00;
mem[16'h8660] = 8'h76;
mem[16'h8661] = 8'h04;
mem[16'h8662] = 8'h03;
mem[16'h8663] = 8'h38;
mem[16'h8664] = 8'h40;
mem[16'h8665] = 8'h03;
mem[16'h8666] = 8'h38;
mem[16'h8667] = 8'h40;
mem[16'h8668] = 8'h03;
mem[16'h8669] = 8'h38;
mem[16'h866A] = 8'h40;
mem[16'h866B] = 8'h03;
mem[16'h866C] = 8'h76;
mem[16'h866D] = 8'h04;
mem[16'h866E] = 8'h03;
mem[16'h866F] = 8'h6E;
mem[16'h8670] = 8'h79;
mem[16'h8671] = 8'h00;
mem[16'h8672] = 8'h00;
mem[16'h8673] = 8'h60;
mem[16'h8674] = 8'h03;
mem[16'h8675] = 8'h00;
mem[16'h8676] = 8'h40;
mem[16'h8677] = 8'h07;
mem[16'h8678] = 8'h5C;
mem[16'h8679] = 8'h73;
mem[16'h867A] = 8'h01;
mem[16'h867B] = 8'h6C;
mem[16'h867C] = 8'h09;
mem[16'h867D] = 8'h06;
mem[16'h867E] = 8'h70;
mem[16'h867F] = 8'h00;
mem[16'h8680] = 8'h07;
mem[16'h8681] = 8'h70;
mem[16'h8682] = 8'h00;
mem[16'h8683] = 8'h07;
mem[16'h8684] = 8'h70;
mem[16'h8685] = 8'h00;
mem[16'h8686] = 8'h07;
mem[16'h8687] = 8'h6C;
mem[16'h8688] = 8'h09;
mem[16'h8689] = 8'h06;
mem[16'h868A] = 8'h5C;
mem[16'h868B] = 8'h73;
mem[16'h868C] = 8'h01;
mem[16'h868D] = 8'h00;
mem[16'h868E] = 8'h40;
mem[16'h868F] = 8'h07;
mem[16'h8690] = 8'h00;
mem[16'h8691] = 8'h00;
mem[16'h8692] = 8'h0F;
mem[16'h8693] = 8'h38;
mem[16'h8694] = 8'h67;
mem[16'h8695] = 8'h03;
mem[16'h8696] = 8'h58;
mem[16'h8697] = 8'h13;
mem[16'h8698] = 8'h0C;
mem[16'h8699] = 8'h60;
mem[16'h869A] = 8'h01;
mem[16'h869B] = 8'h0E;
mem[16'h869C] = 8'h60;
mem[16'h869D] = 8'h01;
mem[16'h869E] = 8'h0E;
mem[16'h869F] = 8'h60;
mem[16'h86A0] = 8'h01;
mem[16'h86A1] = 8'h0E;
mem[16'h86A2] = 8'h58;
mem[16'h86A3] = 8'h13;
mem[16'h86A4] = 8'h0C;
mem[16'h86A5] = 8'h38;
mem[16'h86A6] = 8'h67;
mem[16'h86A7] = 8'h03;
mem[16'h86A8] = 8'h00;
mem[16'h86A9] = 8'h00;
mem[16'h86AA] = 8'h0F;
mem[16'h86AB] = 8'h00;
mem[16'h86AC] = 8'h00;
mem[16'h86AD] = 8'h1E;
mem[16'h86AE] = 8'h70;
mem[16'h86AF] = 8'h4E;
mem[16'h86B0] = 8'h07;
mem[16'h86B1] = 8'h30;
mem[16'h86B2] = 8'h27;
mem[16'h86B3] = 8'h18;
mem[16'h86B4] = 8'h40;
mem[16'h86B5] = 8'h03;
mem[16'h86B6] = 8'h1C;
mem[16'h86B7] = 8'h40;
mem[16'h86B8] = 8'h03;
mem[16'h86B9] = 8'h1C;
mem[16'h86BA] = 8'h40;
mem[16'h86BB] = 8'h03;
mem[16'h86BC] = 8'h1C;
mem[16'h86BD] = 8'h30;
mem[16'h86BE] = 8'h27;
mem[16'h86BF] = 8'h18;
mem[16'h86C0] = 8'h70;
mem[16'h86C1] = 8'h4E;
mem[16'h86C2] = 8'h07;
mem[16'h86C3] = 8'h00;
mem[16'h86C4] = 8'h00;
mem[16'h86C5] = 8'h1E;
mem[16'h86C6] = 8'h00;
mem[16'h86C7] = 8'h00;
mem[16'h86C8] = 8'h3C;
mem[16'h86C9] = 8'h60;
mem[16'h86CA] = 8'h1D;
mem[16'h86CB] = 8'h0F;
mem[16'h86CC] = 8'h60;
mem[16'h86CD] = 8'h4E;
mem[16'h86CE] = 8'h30;
mem[16'h86CF] = 8'h00;
mem[16'h86D0] = 8'h07;
mem[16'h86D1] = 8'h38;
mem[16'h86D2] = 8'h00;
mem[16'h86D3] = 8'h07;
mem[16'h86D4] = 8'h38;
mem[16'h86D5] = 8'h00;
mem[16'h86D6] = 8'h07;
mem[16'h86D7] = 8'h38;
mem[16'h86D8] = 8'h60;
mem[16'h86D9] = 8'h4E;
mem[16'h86DA] = 8'h30;
mem[16'h86DB] = 8'h60;
mem[16'h86DC] = 8'h1D;
mem[16'h86DD] = 8'h0F;
mem[16'h86DE] = 8'h00;
mem[16'h86DF] = 8'h00;
mem[16'h86E0] = 8'h3C;
mem[16'h86E1] = 8'h00;
mem[16'h86E2] = 8'h00;
mem[16'h86E3] = 8'h78;
mem[16'h86E4] = 8'h40;
mem[16'h86E5] = 8'h3B;
mem[16'h86E6] = 8'h1E;
mem[16'h86E7] = 8'h40;
mem[16'h86E8] = 8'h1D;
mem[16'h86E9] = 8'h61;
mem[16'h86EA] = 8'h00;
mem[16'h86EB] = 8'h0E;
mem[16'h86EC] = 8'h70;
mem[16'h86ED] = 8'h00;
mem[16'h86EE] = 8'h0E;
mem[16'h86EF] = 8'h70;
mem[16'h86F0] = 8'h00;
mem[16'h86F1] = 8'h0E;
mem[16'h86F2] = 8'h70;
mem[16'h86F3] = 8'h40;
mem[16'h86F4] = 8'h1D;
mem[16'h86F5] = 8'h61;
mem[16'h86F6] = 8'h40;
mem[16'h86F7] = 8'h3B;
mem[16'h86F8] = 8'h1E;
mem[16'h86F9] = 8'h00;
mem[16'h86FA] = 8'h00;
mem[16'h86FB] = 8'h78;
mem[16'h86FC] = 8'hAD;
mem[16'h86FD] = 8'h14;
mem[16'h86FE] = 8'h87;
mem[16'h86FF] = 8'h29;
mem[16'h8700] = 8'h01;
mem[16'h8701] = 8'h85;
mem[16'h8702] = 8'h60;
mem[16'h8703] = 8'hAD;
mem[16'h8704] = 8'h13;
mem[16'h8705] = 8'h87;
mem[16'h8706] = 8'h6A;
mem[16'h8707] = 8'h29;
mem[16'h8708] = 8'h01;
mem[16'h8709] = 8'h45;
mem[16'h870A] = 8'h60;
mem[16'h870B] = 8'h6A;
mem[16'h870C] = 8'h6E;
mem[16'h870D] = 8'h13;
mem[16'h870E] = 8'h87;
mem[16'h870F] = 8'h6E;
mem[16'h8710] = 8'h14;
mem[16'h8711] = 8'h87;
mem[16'h8712] = 8'h60;
mem[16'h8713] = 8'h5C;
mem[16'h8714] = 8'h9A;
mem[16'h8715] = 8'h00;
mem[16'h8716] = 8'h00;
mem[16'h8717] = 8'h40;
mem[16'h8718] = 8'h02;
mem[16'h8719] = 8'h00;
mem[16'h871A] = 8'h00;
mem[16'h871B] = 8'h00;
mem[16'h871C] = 8'h03;
mem[16'h871D] = 8'h03;
mem[16'h871E] = 8'h00;
mem[16'h871F] = 8'h00;
mem[16'h8720] = 8'h06;
mem[16'h8721] = 8'h00;
mem[16'h8722] = 8'h03;
mem[16'h8723] = 8'h00;
mem[16'h8724] = 8'h03;
mem[16'h8725] = 8'h00;
mem[16'h8726] = 8'h00;
mem[16'h8727] = 8'h03;
mem[16'h8728] = 8'h00;
mem[16'h8729] = 8'h0C;
mem[16'h872A] = 8'h00;
mem[16'h872B] = 8'h00;
mem[16'h872C] = 8'h03;
mem[16'h872D] = 8'h00;
mem[16'h872E] = 8'h00;
mem[16'h872F] = 8'h18;
mem[16'h8730] = 8'h00;
mem[16'h8731] = 8'h03;
mem[16'h8732] = 8'h00;
mem[16'h8733] = 8'h00;
mem[16'h8734] = 8'h00;
mem[16'h8735] = 8'h00;
mem[16'h8736] = 8'h05;
mem[16'h8737] = 8'h00;
mem[16'h8738] = 8'h00;
mem[16'h8739] = 8'h00;
mem[16'h873A] = 8'h06;
mem[16'h873B] = 8'h06;
mem[16'h873C] = 8'h00;
mem[16'h873D] = 8'h00;
mem[16'h873E] = 8'h0C;
mem[16'h873F] = 8'h00;
mem[16'h8740] = 8'h06;
mem[16'h8741] = 8'h00;
mem[16'h8742] = 8'h06;
mem[16'h8743] = 8'h00;
mem[16'h8744] = 8'h00;
mem[16'h8745] = 8'h06;
mem[16'h8746] = 8'h00;
mem[16'h8747] = 8'h18;
mem[16'h8748] = 8'h00;
mem[16'h8749] = 8'h00;
mem[16'h874A] = 8'h06;
mem[16'h874B] = 8'h00;
mem[16'h874C] = 8'h00;
mem[16'h874D] = 8'h30;
mem[16'h874E] = 8'h00;
mem[16'h874F] = 8'h06;
mem[16'h8750] = 8'h00;
mem[16'h8751] = 8'h00;
mem[16'h8752] = 8'h00;
mem[16'h8753] = 8'h00;
mem[16'h8754] = 8'h0A;
mem[16'h8755] = 8'h00;
mem[16'h8756] = 8'h00;
mem[16'h8757] = 8'h00;
mem[16'h8758] = 8'h0C;
mem[16'h8759] = 8'h0C;
mem[16'h875A] = 8'h00;
mem[16'h875B] = 8'h00;
mem[16'h875C] = 8'h18;
mem[16'h875D] = 8'h00;
mem[16'h875E] = 8'h0C;
mem[16'h875F] = 8'h00;
mem[16'h8760] = 8'h0C;
mem[16'h8761] = 8'h00;
mem[16'h8762] = 8'h00;
mem[16'h8763] = 8'h0C;
mem[16'h8764] = 8'h00;
mem[16'h8765] = 8'h30;
mem[16'h8766] = 8'h00;
mem[16'h8767] = 8'h00;
mem[16'h8768] = 8'h0C;
mem[16'h8769] = 8'h00;
mem[16'h876A] = 8'h00;
mem[16'h876B] = 8'h60;
mem[16'h876C] = 8'h00;
mem[16'h876D] = 8'h0C;
mem[16'h876E] = 8'h00;
mem[16'h876F] = 8'h00;
mem[16'h8770] = 8'h00;
mem[16'h8771] = 8'h00;
mem[16'h8772] = 8'h14;
mem[16'h8773] = 8'h00;
mem[16'h8774] = 8'h00;
mem[16'h8775] = 8'h00;
mem[16'h8776] = 8'h18;
mem[16'h8777] = 8'h18;
mem[16'h8778] = 8'h00;
mem[16'h8779] = 8'h00;
mem[16'h877A] = 8'h30;
mem[16'h877B] = 8'h00;
mem[16'h877C] = 8'h18;
mem[16'h877D] = 8'h00;
mem[16'h877E] = 8'h18;
mem[16'h877F] = 8'h00;
mem[16'h8780] = 8'h00;
mem[16'h8781] = 8'h18;
mem[16'h8782] = 8'h00;
mem[16'h8783] = 8'h60;
mem[16'h8784] = 8'h00;
mem[16'h8785] = 8'h00;
mem[16'h8786] = 8'h18;
mem[16'h8787] = 8'h00;
mem[16'h8788] = 8'h00;
mem[16'h8789] = 8'h40;
mem[16'h878A] = 8'h01;
mem[16'h878B] = 8'h18;
mem[16'h878C] = 8'h00;
mem[16'h878D] = 8'h00;
mem[16'h878E] = 8'h00;
mem[16'h878F] = 8'h00;
mem[16'h8790] = 8'h28;
mem[16'h8791] = 8'h00;
mem[16'h8792] = 8'h00;
mem[16'h8793] = 8'h00;
mem[16'h8794] = 8'h30;
mem[16'h8795] = 8'h30;
mem[16'h8796] = 8'h00;
mem[16'h8797] = 8'h00;
mem[16'h8798] = 8'h60;
mem[16'h8799] = 8'h00;
mem[16'h879A] = 8'h30;
mem[16'h879B] = 8'h00;
mem[16'h879C] = 8'h30;
mem[16'h879D] = 8'h00;
mem[16'h879E] = 8'h00;
mem[16'h879F] = 8'h30;
mem[16'h87A0] = 8'h00;
mem[16'h87A1] = 8'h40;
mem[16'h87A2] = 8'h01;
mem[16'h87A3] = 8'h00;
mem[16'h87A4] = 8'h30;
mem[16'h87A5] = 8'h00;
mem[16'h87A6] = 8'h00;
mem[16'h87A7] = 8'h00;
mem[16'h87A8] = 8'h03;
mem[16'h87A9] = 8'h30;
mem[16'h87AA] = 8'h00;
mem[16'h87AB] = 8'h00;
mem[16'h87AC] = 8'h00;
mem[16'h87AD] = 8'h00;
mem[16'h87AE] = 8'h50;
mem[16'h87AF] = 8'h00;
mem[16'h87B0] = 8'h00;
mem[16'h87B1] = 8'h00;
mem[16'h87B2] = 8'h60;
mem[16'h87B3] = 8'h60;
mem[16'h87B4] = 8'h00;
mem[16'h87B5] = 8'h00;
mem[16'h87B6] = 8'h40;
mem[16'h87B7] = 8'h01;
mem[16'h87B8] = 8'h60;
mem[16'h87B9] = 8'h00;
mem[16'h87BA] = 8'h60;
mem[16'h87BB] = 8'h00;
mem[16'h87BC] = 8'h00;
mem[16'h87BD] = 8'h60;
mem[16'h87BE] = 8'h00;
mem[16'h87BF] = 8'h00;
mem[16'h87C0] = 8'h03;
mem[16'h87C1] = 8'h00;
mem[16'h87C2] = 8'h60;
mem[16'h87C3] = 8'h00;
mem[16'h87C4] = 8'h00;
mem[16'h87C5] = 8'h00;
mem[16'h87C6] = 8'h06;
mem[16'h87C7] = 8'h60;
mem[16'h87C8] = 8'h00;
mem[16'h87C9] = 8'h00;
mem[16'h87CA] = 8'h00;
mem[16'h87CB] = 8'h00;
mem[16'h87CC] = 8'h20;
mem[16'h87CD] = 8'h01;
mem[16'h87CE] = 8'h00;
mem[16'h87CF] = 8'h00;
mem[16'h87D0] = 8'h40;
mem[16'h87D1] = 8'h41;
mem[16'h87D2] = 8'h01;
mem[16'h87D3] = 8'h00;
mem[16'h87D4] = 8'h00;
mem[16'h87D5] = 8'h03;
mem[16'h87D6] = 8'h40;
mem[16'h87D7] = 8'h01;
mem[16'h87D8] = 8'h40;
mem[16'h87D9] = 8'h01;
mem[16'h87DA] = 8'h00;
mem[16'h87DB] = 8'h40;
mem[16'h87DC] = 8'h01;
mem[16'h87DD] = 8'h00;
mem[16'h87DE] = 8'h06;
mem[16'h87DF] = 8'h00;
mem[16'h87E0] = 8'h40;
mem[16'h87E1] = 8'h01;
mem[16'h87E2] = 8'h00;
mem[16'h87E3] = 8'h00;
mem[16'h87E4] = 8'h0C;
mem[16'h87E5] = 8'h40;
mem[16'h87E6] = 8'h01;
mem[16'h87E7] = 8'h00;
mem[16'h87E8] = 8'h00;
mem[16'h87E9] = 8'h58;
mem[16'h87EA] = 8'h01;
mem[16'h87EB] = 8'h00;
mem[16'h87EC] = 8'h40;
mem[16'h87ED] = 8'h41;
mem[16'h87EE] = 8'h01;
mem[16'h87EF] = 8'h40;
mem[16'h87F0] = 8'h01;
mem[16'h87F1] = 8'h40;
mem[16'h87F2] = 8'h01;
mem[16'h87F3] = 8'h40;
mem[16'h87F4] = 8'h01;
mem[16'h87F5] = 8'h40;
mem[16'h87F6] = 8'h01;
mem[16'h87F7] = 8'h40;
mem[16'h87F8] = 8'h01;
mem[16'h87F9] = 8'h40;
mem[16'h87FA] = 8'h01;
mem[16'h87FB] = 8'h40;
mem[16'h87FC] = 8'h01;
mem[16'h87FD] = 8'h40;
mem[16'h87FE] = 8'h01;
mem[16'h87FF] = 8'h40;
mem[16'h8800] = 8'h01;
mem[16'h8801] = 8'h40;
mem[16'h8802] = 8'h01;
mem[16'h8803] = 8'h40;
mem[16'h8804] = 8'h01;
mem[16'h8805] = 8'h40;
mem[16'h8806] = 8'h01;
mem[16'h8807] = 8'h00;
mem[16'h8808] = 8'h00;
mem[16'h8809] = 8'h6C;
mem[16'h880A] = 8'h00;
mem[16'h880B] = 8'h00;
mem[16'h880C] = 8'h60;
mem[16'h880D] = 8'h60;
mem[16'h880E] = 8'h00;
mem[16'h880F] = 8'h60;
mem[16'h8810] = 8'h00;
mem[16'h8811] = 8'h60;
mem[16'h8812] = 8'h00;
mem[16'h8813] = 8'h60;
mem[16'h8814] = 8'h00;
mem[16'h8815] = 8'h60;
mem[16'h8816] = 8'h00;
mem[16'h8817] = 8'h60;
mem[16'h8818] = 8'h00;
mem[16'h8819] = 8'h60;
mem[16'h881A] = 8'h00;
mem[16'h881B] = 8'h60;
mem[16'h881C] = 8'h00;
mem[16'h881D] = 8'h60;
mem[16'h881E] = 8'h00;
mem[16'h881F] = 8'h60;
mem[16'h8820] = 8'h00;
mem[16'h8821] = 8'h60;
mem[16'h8822] = 8'h00;
mem[16'h8823] = 8'h60;
mem[16'h8824] = 8'h00;
mem[16'h8825] = 8'h60;
mem[16'h8826] = 8'h00;
mem[16'h8827] = 8'h00;
mem[16'h8828] = 8'h00;
mem[16'h8829] = 8'h36;
mem[16'h882A] = 8'h00;
mem[16'h882B] = 8'h00;
mem[16'h882C] = 8'h30;
mem[16'h882D] = 8'h30;
mem[16'h882E] = 8'h00;
mem[16'h882F] = 8'h30;
mem[16'h8830] = 8'h00;
mem[16'h8831] = 8'h30;
mem[16'h8832] = 8'h00;
mem[16'h8833] = 8'h30;
mem[16'h8834] = 8'h00;
mem[16'h8835] = 8'h30;
mem[16'h8836] = 8'h00;
mem[16'h8837] = 8'h30;
mem[16'h8838] = 8'h00;
mem[16'h8839] = 8'h30;
mem[16'h883A] = 8'h00;
mem[16'h883B] = 8'h30;
mem[16'h883C] = 8'h00;
mem[16'h883D] = 8'h30;
mem[16'h883E] = 8'h00;
mem[16'h883F] = 8'h30;
mem[16'h8840] = 8'h00;
mem[16'h8841] = 8'h30;
mem[16'h8842] = 8'h00;
mem[16'h8843] = 8'h30;
mem[16'h8844] = 8'h00;
mem[16'h8845] = 8'h30;
mem[16'h8846] = 8'h00;
mem[16'h8847] = 8'h00;
mem[16'h8848] = 8'h00;
mem[16'h8849] = 8'h1B;
mem[16'h884A] = 8'h00;
mem[16'h884B] = 8'h00;
mem[16'h884C] = 8'h18;
mem[16'h884D] = 8'h18;
mem[16'h884E] = 8'h00;
mem[16'h884F] = 8'h18;
mem[16'h8850] = 8'h00;
mem[16'h8851] = 8'h18;
mem[16'h8852] = 8'h00;
mem[16'h8853] = 8'h18;
mem[16'h8854] = 8'h00;
mem[16'h8855] = 8'h18;
mem[16'h8856] = 8'h00;
mem[16'h8857] = 8'h18;
mem[16'h8858] = 8'h00;
mem[16'h8859] = 8'h18;
mem[16'h885A] = 8'h00;
mem[16'h885B] = 8'h18;
mem[16'h885C] = 8'h00;
mem[16'h885D] = 8'h18;
mem[16'h885E] = 8'h00;
mem[16'h885F] = 8'h18;
mem[16'h8860] = 8'h00;
mem[16'h8861] = 8'h18;
mem[16'h8862] = 8'h00;
mem[16'h8863] = 8'h18;
mem[16'h8864] = 8'h00;
mem[16'h8865] = 8'h18;
mem[16'h8866] = 8'h00;
mem[16'h8867] = 8'h00;
mem[16'h8868] = 8'h40;
mem[16'h8869] = 8'h0D;
mem[16'h886A] = 8'h00;
mem[16'h886B] = 8'h00;
mem[16'h886C] = 8'h0C;
mem[16'h886D] = 8'h0C;
mem[16'h886E] = 8'h00;
mem[16'h886F] = 8'h0C;
mem[16'h8870] = 8'h00;
mem[16'h8871] = 8'h0C;
mem[16'h8872] = 8'h00;
mem[16'h8873] = 8'h0C;
mem[16'h8874] = 8'h00;
mem[16'h8875] = 8'h0C;
mem[16'h8876] = 8'h00;
mem[16'h8877] = 8'h0C;
mem[16'h8878] = 8'h00;
mem[16'h8879] = 8'h0C;
mem[16'h887A] = 8'h00;
mem[16'h887B] = 8'h0C;
mem[16'h887C] = 8'h00;
mem[16'h887D] = 8'h0C;
mem[16'h887E] = 8'h00;
mem[16'h887F] = 8'h0C;
mem[16'h8880] = 8'h00;
mem[16'h8881] = 8'h0C;
mem[16'h8882] = 8'h00;
mem[16'h8883] = 8'h0C;
mem[16'h8884] = 8'h00;
mem[16'h8885] = 8'h0C;
mem[16'h8886] = 8'h00;
mem[16'h8887] = 8'h00;
mem[16'h8888] = 8'h60;
mem[16'h8889] = 8'h06;
mem[16'h888A] = 8'h00;
mem[16'h888B] = 8'h00;
mem[16'h888C] = 8'h06;
mem[16'h888D] = 8'h06;
mem[16'h888E] = 8'h00;
mem[16'h888F] = 8'h06;
mem[16'h8890] = 8'h00;
mem[16'h8891] = 8'h06;
mem[16'h8892] = 8'h00;
mem[16'h8893] = 8'h06;
mem[16'h8894] = 8'h00;
mem[16'h8895] = 8'h06;
mem[16'h8896] = 8'h00;
mem[16'h8897] = 8'h06;
mem[16'h8898] = 8'h00;
mem[16'h8899] = 8'h06;
mem[16'h889A] = 8'h00;
mem[16'h889B] = 8'h06;
mem[16'h889C] = 8'h00;
mem[16'h889D] = 8'h06;
mem[16'h889E] = 8'h00;
mem[16'h889F] = 8'h06;
mem[16'h88A0] = 8'h00;
mem[16'h88A1] = 8'h06;
mem[16'h88A2] = 8'h00;
mem[16'h88A3] = 8'h06;
mem[16'h88A4] = 8'h00;
mem[16'h88A5] = 8'h06;
mem[16'h88A6] = 8'h00;
mem[16'h88A7] = 8'h00;
mem[16'h88A8] = 8'h30;
mem[16'h88A9] = 8'h03;
mem[16'h88AA] = 8'h00;
mem[16'h88AB] = 8'h00;
mem[16'h88AC] = 8'h03;
mem[16'h88AD] = 8'h03;
mem[16'h88AE] = 8'h00;
mem[16'h88AF] = 8'h03;
mem[16'h88B0] = 8'h00;
mem[16'h88B1] = 8'h03;
mem[16'h88B2] = 8'h00;
mem[16'h88B3] = 8'h03;
mem[16'h88B4] = 8'h00;
mem[16'h88B5] = 8'h03;
mem[16'h88B6] = 8'h00;
mem[16'h88B7] = 8'h03;
mem[16'h88B8] = 8'h00;
mem[16'h88B9] = 8'h03;
mem[16'h88BA] = 8'h00;
mem[16'h88BB] = 8'h03;
mem[16'h88BC] = 8'h00;
mem[16'h88BD] = 8'h03;
mem[16'h88BE] = 8'h00;
mem[16'h88BF] = 8'h03;
mem[16'h88C0] = 8'h00;
mem[16'h88C1] = 8'h03;
mem[16'h88C2] = 8'h00;
mem[16'h88C3] = 8'h03;
mem[16'h88C4] = 8'h00;
mem[16'h88C5] = 8'h03;
mem[16'h88C6] = 8'h00;
mem[16'h88C7] = 8'h00;
mem[16'h88C8] = 8'h00;
mem[16'h88C9] = 8'h28;
mem[16'h88CA] = 8'h00;
mem[16'h88CB] = 8'h00;
mem[16'h88CC] = 8'h36;
mem[16'h88CD] = 8'h40;
mem[16'h88CE] = 8'h47;
mem[16'h88CF] = 8'h25;
mem[16'h88D0] = 8'h40;
mem[16'h88D1] = 8'h01;
mem[16'h88D2] = 8'h24;
mem[16'h88D3] = 8'h40;
mem[16'h88D4] = 8'h04;
mem[16'h88D5] = 8'h09;
mem[16'h88D6] = 8'h40;
mem[16'h88D7] = 8'h61;
mem[16'h88D8] = 8'h0A;
mem[16'h88D9] = 8'h40;
mem[16'h88DA] = 8'h59;
mem[16'h88DB] = 8'h2A;
mem[16'h88DC] = 8'h40;
mem[16'h88DD] = 8'h53;
mem[16'h88DE] = 8'h2A;
mem[16'h88DF] = 8'h40;
mem[16'h88E0] = 8'h01;
mem[16'h88E1] = 8'h30;
mem[16'h88E2] = 8'h40;
mem[16'h88E3] = 8'h01;
mem[16'h88E4] = 8'h0C;
mem[16'h88E5] = 8'h00;
mem[16'h88E6] = 8'h00;
mem[16'h88E7] = 8'h14;
mem[16'h88E8] = 8'h00;
mem[16'h88E9] = 8'h00;
mem[16'h88EA] = 8'h1B;
mem[16'h88EB] = 8'h60;
mem[16'h88EC] = 8'h63;
mem[16'h88ED] = 8'h12;
mem[16'h88EE] = 8'h60;
mem[16'h88EF] = 8'h00;
mem[16'h88F0] = 8'h12;
mem[16'h88F1] = 8'h20;
mem[16'h88F2] = 8'h42;
mem[16'h88F3] = 8'h04;
mem[16'h88F4] = 8'h60;
mem[16'h88F5] = 8'h30;
mem[16'h88F6] = 8'h05;
mem[16'h88F7] = 8'h60;
mem[16'h88F8] = 8'h2C;
mem[16'h88F9] = 8'h15;
mem[16'h88FA] = 8'h60;
mem[16'h88FB] = 8'h29;
mem[16'h88FC] = 8'h15;
mem[16'h88FD] = 8'h60;
mem[16'h88FE] = 8'h00;
mem[16'h88FF] = 8'h18;
mem[16'h8900] = 8'h60;
mem[16'h8901] = 8'h00;
mem[16'h8902] = 8'h06;
mem[16'h8903] = 8'h00;
mem[16'h8904] = 8'h00;
mem[16'h8905] = 8'h0A;
mem[16'h8906] = 8'h00;
mem[16'h8907] = 8'h40;
mem[16'h8908] = 8'h0D;
mem[16'h8909] = 8'h70;
mem[16'h890A] = 8'h31;
mem[16'h890B] = 8'h09;
mem[16'h890C] = 8'h30;
mem[16'h890D] = 8'h00;
mem[16'h890E] = 8'h09;
mem[16'h890F] = 8'h10;
mem[16'h8910] = 8'h21;
mem[16'h8911] = 8'h02;
mem[16'h8912] = 8'h30;
mem[16'h8913] = 8'h58;
mem[16'h8914] = 8'h02;
mem[16'h8915] = 8'h30;
mem[16'h8916] = 8'h56;
mem[16'h8917] = 8'h0A;
mem[16'h8918] = 8'h70;
mem[16'h8919] = 8'h54;
mem[16'h891A] = 8'h0A;
mem[16'h891B] = 8'h30;
mem[16'h891C] = 8'h00;
mem[16'h891D] = 8'h0C;
mem[16'h891E] = 8'h30;
mem[16'h891F] = 8'h00;
mem[16'h8920] = 8'h03;
mem[16'h8921] = 8'h00;
mem[16'h8922] = 8'h00;
mem[16'h8923] = 8'h05;
mem[16'h8924] = 8'h00;
mem[16'h8925] = 8'h60;
mem[16'h8926] = 8'h06;
mem[16'h8927] = 8'h78;
mem[16'h8928] = 8'h58;
mem[16'h8929] = 8'h04;
mem[16'h892A] = 8'h18;
mem[16'h892B] = 8'h40;
mem[16'h892C] = 8'h04;
mem[16'h892D] = 8'h48;
mem[16'h892E] = 8'h10;
mem[16'h892F] = 8'h01;
mem[16'h8930] = 8'h18;
mem[16'h8931] = 8'h2C;
mem[16'h8932] = 8'h01;
mem[16'h8933] = 8'h18;
mem[16'h8934] = 8'h2B;
mem[16'h8935] = 8'h05;
mem[16'h8936] = 8'h38;
mem[16'h8937] = 8'h2A;
mem[16'h8938] = 8'h05;
mem[16'h8939] = 8'h18;
mem[16'h893A] = 8'h00;
mem[16'h893B] = 8'h06;
mem[16'h893C] = 8'h18;
mem[16'h893D] = 8'h40;
mem[16'h893E] = 8'h01;
mem[16'h893F] = 8'h00;
mem[16'h8940] = 8'h40;
mem[16'h8941] = 8'h02;
mem[16'h8942] = 8'h00;
mem[16'h8943] = 8'h30;
mem[16'h8944] = 8'h03;
mem[16'h8945] = 8'h3C;
mem[16'h8946] = 8'h2C;
mem[16'h8947] = 8'h02;
mem[16'h8948] = 8'h0C;
mem[16'h8949] = 8'h20;
mem[16'h894A] = 8'h02;
mem[16'h894B] = 8'h24;
mem[16'h894C] = 8'h48;
mem[16'h894D] = 8'h00;
mem[16'h894E] = 8'h0C;
mem[16'h894F] = 8'h56;
mem[16'h8950] = 8'h00;
mem[16'h8951] = 8'h4C;
mem[16'h8952] = 8'h55;
mem[16'h8953] = 8'h02;
mem[16'h8954] = 8'h1C;
mem[16'h8955] = 8'h55;
mem[16'h8956] = 8'h02;
mem[16'h8957] = 8'h0C;
mem[16'h8958] = 8'h00;
mem[16'h8959] = 8'h03;
mem[16'h895A] = 8'h0C;
mem[16'h895B] = 8'h60;
mem[16'h895C] = 8'h00;
mem[16'h895D] = 8'h00;
mem[16'h895E] = 8'h20;
mem[16'h895F] = 8'h01;
mem[16'h8960] = 8'h00;
mem[16'h8961] = 8'h58;
mem[16'h8962] = 8'h01;
mem[16'h8963] = 8'h1E;
mem[16'h8964] = 8'h16;
mem[16'h8965] = 8'h01;
mem[16'h8966] = 8'h06;
mem[16'h8967] = 8'h10;
mem[16'h8968] = 8'h01;
mem[16'h8969] = 8'h12;
mem[16'h896A] = 8'h24;
mem[16'h896B] = 8'h00;
mem[16'h896C] = 8'h06;
mem[16'h896D] = 8'h2B;
mem[16'h896E] = 8'h00;
mem[16'h896F] = 8'h66;
mem[16'h8970] = 8'h2A;
mem[16'h8971] = 8'h01;
mem[16'h8972] = 8'h4E;
mem[16'h8973] = 8'h2A;
mem[16'h8974] = 8'h01;
mem[16'h8975] = 8'h06;
mem[16'h8976] = 8'h40;
mem[16'h8977] = 8'h01;
mem[16'h8978] = 8'h06;
mem[16'h8979] = 8'h30;
mem[16'h897A] = 8'h00;
mem[16'h897B] = 8'h00;
mem[16'h897C] = 8'h50;
mem[16'h897D] = 8'h00;
mem[16'h897E] = 8'h00;
mem[16'h897F] = 8'h6C;
mem[16'h8980] = 8'h00;
mem[16'h8981] = 8'h0F;
mem[16'h8982] = 8'h4B;
mem[16'h8983] = 8'h00;
mem[16'h8984] = 8'h03;
mem[16'h8985] = 8'h48;
mem[16'h8986] = 8'h00;
mem[16'h8987] = 8'h09;
mem[16'h8988] = 8'h12;
mem[16'h8989] = 8'h00;
mem[16'h898A] = 8'h43;
mem[16'h898B] = 8'h15;
mem[16'h898C] = 8'h00;
mem[16'h898D] = 8'h33;
mem[16'h898E] = 8'h55;
mem[16'h898F] = 8'h00;
mem[16'h8990] = 8'h27;
mem[16'h8991] = 8'h55;
mem[16'h8992] = 8'h00;
mem[16'h8993] = 8'h03;
mem[16'h8994] = 8'h60;
mem[16'h8995] = 8'h00;
mem[16'h8996] = 8'h03;
mem[16'h8997] = 8'h18;
mem[16'h8998] = 8'h00;
mem[16'h8999] = 8'h40;
mem[16'h899A] = 8'h07;
mem[16'h899B] = 8'h00;
mem[16'h899C] = 8'h00;
mem[16'h899D] = 8'h40;
mem[16'h899E] = 8'h19;
mem[16'h899F] = 8'h00;
mem[16'h89A0] = 8'h00;
mem[16'h89A1] = 8'h40;
mem[16'h89A2] = 8'h1C;
mem[16'h89A3] = 8'h00;
mem[16'h89A4] = 8'h00;
mem[16'h89A5] = 8'h40;
mem[16'h89A6] = 8'h61;
mem[16'h89A7] = 8'h00;
mem[16'h89A8] = 8'h00;
mem[16'h89A9] = 8'h40;
mem[16'h89AA] = 8'h01;
mem[16'h89AB] = 8'h40;
mem[16'h89AC] = 8'h01;
mem[16'h89AD] = 8'h40;
mem[16'h89AE] = 8'h09;
mem[16'h89AF] = 8'h00;
mem[16'h89B0] = 8'h01;
mem[16'h89B1] = 8'h40;
mem[16'h89B2] = 8'h01;
mem[16'h89B3] = 8'h40;
mem[16'h89B4] = 8'h01;
mem[16'h89B5] = 8'h40;
mem[16'h89B6] = 8'h01;
mem[16'h89B7] = 8'h30;
mem[16'h89B8] = 8'h00;
mem[16'h89B9] = 8'h60;
mem[16'h89BA] = 8'h03;
mem[16'h89BB] = 8'h00;
mem[16'h89BC] = 8'h00;
mem[16'h89BD] = 8'h60;
mem[16'h89BE] = 8'h0C;
mem[16'h89BF] = 8'h00;
mem[16'h89C0] = 8'h00;
mem[16'h89C1] = 8'h20;
mem[16'h89C2] = 8'h0E;
mem[16'h89C3] = 8'h00;
mem[16'h89C4] = 8'h00;
mem[16'h89C5] = 8'h60;
mem[16'h89C6] = 8'h30;
mem[16'h89C7] = 8'h00;
mem[16'h89C8] = 8'h00;
mem[16'h89C9] = 8'h60;
mem[16'h89CA] = 8'h00;
mem[16'h89CB] = 8'h60;
mem[16'h89CC] = 8'h00;
mem[16'h89CD] = 8'h60;
mem[16'h89CE] = 8'h04;
mem[16'h89CF] = 8'h40;
mem[16'h89D0] = 8'h00;
mem[16'h89D1] = 8'h60;
mem[16'h89D2] = 8'h00;
mem[16'h89D3] = 8'h60;
mem[16'h89D4] = 8'h00;
mem[16'h89D5] = 8'h60;
mem[16'h89D6] = 8'h00;
mem[16'h89D7] = 8'h18;
mem[16'h89D8] = 8'h00;
mem[16'h89D9] = 8'h70;
mem[16'h89DA] = 8'h01;
mem[16'h89DB] = 8'h00;
mem[16'h89DC] = 8'h00;
mem[16'h89DD] = 8'h30;
mem[16'h89DE] = 8'h06;
mem[16'h89DF] = 8'h00;
mem[16'h89E0] = 8'h00;
mem[16'h89E1] = 8'h10;
mem[16'h89E2] = 8'h07;
mem[16'h89E3] = 8'h00;
mem[16'h89E4] = 8'h00;
mem[16'h89E5] = 8'h30;
mem[16'h89E6] = 8'h18;
mem[16'h89E7] = 8'h00;
mem[16'h89E8] = 8'h00;
mem[16'h89E9] = 8'h30;
mem[16'h89EA] = 8'h00;
mem[16'h89EB] = 8'h30;
mem[16'h89EC] = 8'h00;
mem[16'h89ED] = 8'h30;
mem[16'h89EE] = 8'h02;
mem[16'h89EF] = 8'h20;
mem[16'h89F0] = 8'h00;
mem[16'h89F1] = 8'h30;
mem[16'h89F2] = 8'h00;
mem[16'h89F3] = 8'h30;
mem[16'h89F4] = 8'h00;
mem[16'h89F5] = 8'h30;
mem[16'h89F6] = 8'h00;
mem[16'h89F7] = 8'h0C;
mem[16'h89F8] = 8'h00;
mem[16'h89F9] = 8'h78;
mem[16'h89FA] = 8'h00;
mem[16'h89FB] = 8'h00;
mem[16'h89FC] = 8'h00;
mem[16'h89FD] = 8'h18;
mem[16'h89FE] = 8'h03;
mem[16'h89FF] = 8'h00;
mem[16'h8A00] = 8'h00;
mem[16'h8A01] = 8'h48;
mem[16'h8A02] = 8'h03;
mem[16'h8A03] = 8'h00;
mem[16'h8A04] = 8'h00;
mem[16'h8A05] = 8'h18;
mem[16'h8A06] = 8'h0C;
mem[16'h8A07] = 8'h00;
mem[16'h8A08] = 8'h00;
mem[16'h8A09] = 8'h18;
mem[16'h8A0A] = 8'h00;
mem[16'h8A0B] = 8'h18;
mem[16'h8A0C] = 8'h00;
mem[16'h8A0D] = 8'h18;
mem[16'h8A0E] = 8'h01;
mem[16'h8A0F] = 8'h10;
mem[16'h8A10] = 8'h00;
mem[16'h8A11] = 8'h18;
mem[16'h8A12] = 8'h00;
mem[16'h8A13] = 8'h18;
mem[16'h8A14] = 8'h00;
mem[16'h8A15] = 8'h18;
mem[16'h8A16] = 8'h00;
mem[16'h8A17] = 8'h06;
mem[16'h8A18] = 8'h00;
mem[16'h8A19] = 8'h3C;
mem[16'h8A1A] = 8'h00;
mem[16'h8A1B] = 8'h00;
mem[16'h8A1C] = 8'h00;
mem[16'h8A1D] = 8'h4C;
mem[16'h8A1E] = 8'h01;
mem[16'h8A1F] = 8'h00;
mem[16'h8A20] = 8'h00;
mem[16'h8A21] = 8'h64;
mem[16'h8A22] = 8'h01;
mem[16'h8A23] = 8'h00;
mem[16'h8A24] = 8'h00;
mem[16'h8A25] = 8'h0C;
mem[16'h8A26] = 8'h06;
mem[16'h8A27] = 8'h00;
mem[16'h8A28] = 8'h00;
mem[16'h8A29] = 8'h0C;
mem[16'h8A2A] = 8'h00;
mem[16'h8A2B] = 8'h0C;
mem[16'h8A2C] = 8'h00;
mem[16'h8A2D] = 8'h4C;
mem[16'h8A2E] = 8'h00;
mem[16'h8A2F] = 8'h08;
mem[16'h8A30] = 8'h00;
mem[16'h8A31] = 8'h0C;
mem[16'h8A32] = 8'h00;
mem[16'h8A33] = 8'h0C;
mem[16'h8A34] = 8'h00;
mem[16'h8A35] = 8'h0C;
mem[16'h8A36] = 8'h00;
mem[16'h8A37] = 8'h03;
mem[16'h8A38] = 8'h00;
mem[16'h8A39] = 8'h1E;
mem[16'h8A3A] = 8'h00;
mem[16'h8A3B] = 8'h00;
mem[16'h8A3C] = 8'h00;
mem[16'h8A3D] = 8'h66;
mem[16'h8A3E] = 8'h00;
mem[16'h8A3F] = 8'h00;
mem[16'h8A40] = 8'h00;
mem[16'h8A41] = 8'h72;
mem[16'h8A42] = 8'h00;
mem[16'h8A43] = 8'h00;
mem[16'h8A44] = 8'h00;
mem[16'h8A45] = 8'h06;
mem[16'h8A46] = 8'h03;
mem[16'h8A47] = 8'h00;
mem[16'h8A48] = 8'h00;
mem[16'h8A49] = 8'h06;
mem[16'h8A4A] = 8'h00;
mem[16'h8A4B] = 8'h06;
mem[16'h8A4C] = 8'h00;
mem[16'h8A4D] = 8'h26;
mem[16'h8A4E] = 8'h00;
mem[16'h8A4F] = 8'h04;
mem[16'h8A50] = 8'h00;
mem[16'h8A51] = 8'h06;
mem[16'h8A52] = 8'h00;
mem[16'h8A53] = 8'h06;
mem[16'h8A54] = 8'h00;
mem[16'h8A55] = 8'h06;
mem[16'h8A56] = 8'h40;
mem[16'h8A57] = 8'h01;
mem[16'h8A58] = 8'h00;
mem[16'h8A59] = 8'h0F;
mem[16'h8A5A] = 8'h00;
mem[16'h8A5B] = 8'h00;
mem[16'h8A5C] = 8'h00;
mem[16'h8A5D] = 8'h33;
mem[16'h8A5E] = 8'h00;
mem[16'h8A5F] = 8'h00;
mem[16'h8A60] = 8'h00;
mem[16'h8A61] = 8'h39;
mem[16'h8A62] = 8'h00;
mem[16'h8A63] = 8'h00;
mem[16'h8A64] = 8'h00;
mem[16'h8A65] = 8'h43;
mem[16'h8A66] = 8'h01;
mem[16'h8A67] = 8'h00;
mem[16'h8A68] = 8'h00;
mem[16'h8A69] = 8'h03;
mem[16'h8A6A] = 8'h00;
mem[16'h8A6B] = 8'h03;
mem[16'h8A6C] = 8'h00;
mem[16'h8A6D] = 8'h13;
mem[16'h8A6E] = 8'h00;
mem[16'h8A6F] = 8'h02;
mem[16'h8A70] = 8'h00;
mem[16'h8A71] = 8'h03;
mem[16'h8A72] = 8'h00;
mem[16'h8A73] = 8'h03;
mem[16'h8A74] = 8'h00;
mem[16'h8A75] = 8'h03;
mem[16'h8A76] = 8'h60;
mem[16'h8A77] = 8'h00;
mem[16'h8A78] = 8'h00;
mem[16'h8A79] = 8'hA2;
mem[16'h8A7A] = 8'h00;
mem[16'h8A7B] = 8'hA4;
mem[16'h8A7C] = 8'h56;
mem[16'h8A7D] = 8'hB9;
mem[16'h8A7E] = 8'hD5;
mem[16'h8A7F] = 8'h8E;
mem[16'h8A80] = 8'h85;
mem[16'h8A81] = 8'h59;
mem[16'h8A82] = 8'hB9;
mem[16'h8A83] = 8'h95;
mem[16'h8A84] = 8'h8F;
mem[16'h8A85] = 8'h85;
mem[16'h8A86] = 8'h5A;
mem[16'h8A87] = 8'hA4;
mem[16'h8A88] = 8'h57;
mem[16'h8A89] = 8'hB9;
mem[16'h8A8A] = 8'h56;
mem[16'h8A8B] = 8'h8D;
mem[16'h8A8C] = 8'hA8;
mem[16'h8A8D] = 8'hBD;
mem[16'h8A8E] = 8'h00;
mem[16'h8A8F] = 8'h00;
mem[16'h8A90] = 8'h29;
mem[16'h8A91] = 8'h80;
mem[16'h8A92] = 8'h85;
mem[16'h8A93] = 8'h6D;
mem[16'h8A94] = 8'hBD;
mem[16'h8A95] = 8'h00;
mem[16'h8A96] = 8'h00;
mem[16'h8A97] = 8'h29;
mem[16'h8A98] = 8'h7F;
mem[16'h8A99] = 8'h51;
mem[16'h8A9A] = 8'h59;
mem[16'h8A9B] = 8'h05;
mem[16'h8A9C] = 8'h6D;
mem[16'h8A9D] = 8'h91;
mem[16'h8A9E] = 8'h59;
mem[16'h8A9F] = 8'hE8;
mem[16'h8AA0] = 8'hC8;
mem[16'h8AA1] = 8'hBD;
mem[16'h8AA2] = 8'h00;
mem[16'h8AA3] = 8'h00;
mem[16'h8AA4] = 8'h29;
mem[16'h8AA5] = 8'h7F;
mem[16'h8AA6] = 8'h51;
mem[16'h8AA7] = 8'h59;
mem[16'h8AA8] = 8'h05;
mem[16'h8AA9] = 8'h6D;
mem[16'h8AAA] = 8'h91;
mem[16'h8AAB] = 8'h59;
mem[16'h8AAC] = 8'hC8;
mem[16'h8AAD] = 8'hE8;
mem[16'h8AAE] = 8'hBD;
mem[16'h8AAF] = 8'h00;
mem[16'h8AB0] = 8'h00;
mem[16'h8AB1] = 8'h29;
mem[16'h8AB2] = 8'h7F;
mem[16'h8AB3] = 8'h51;
mem[16'h8AB4] = 8'h59;
mem[16'h8AB5] = 8'h05;
mem[16'h8AB6] = 8'h6D;
mem[16'h8AB7] = 8'h91;
mem[16'h8AB8] = 8'h59;
mem[16'h8AB9] = 8'hC8;
mem[16'h8ABA] = 8'hE8;
mem[16'h8ABB] = 8'hBD;
mem[16'h8ABC] = 8'h00;
mem[16'h8ABD] = 8'h00;
mem[16'h8ABE] = 8'h29;
mem[16'h8ABF] = 8'h7F;
mem[16'h8AC0] = 8'h51;
mem[16'h8AC1] = 8'h59;
mem[16'h8AC2] = 8'h05;
mem[16'h8AC3] = 8'h6D;
mem[16'h8AC4] = 8'h91;
mem[16'h8AC5] = 8'h59;
mem[16'h8AC6] = 8'hE6;
mem[16'h8AC7] = 8'h56;
mem[16'h8AC8] = 8'hE8;
mem[16'h8AC9] = 8'hE0;
mem[16'h8ACA] = 8'h1E;
mem[16'h8ACB] = 8'hB0;
mem[16'h8ACC] = 8'h03;
mem[16'h8ACD] = 8'h4C;
mem[16'h8ACE] = 8'h7B;
mem[16'h8ACF] = 8'h8A;
mem[16'h8AD0] = 8'h60;
mem[16'h8AD1] = 8'h8D;
mem[16'h8AD2] = 8'h8E;
mem[16'h8AD3] = 8'h8A;
mem[16'h8AD4] = 8'h8D;
mem[16'h8AD5] = 8'h95;
mem[16'h8AD6] = 8'h8A;
mem[16'h8AD7] = 8'h8D;
mem[16'h8AD8] = 8'hA2;
mem[16'h8AD9] = 8'h8A;
mem[16'h8ADA] = 8'h8D;
mem[16'h8ADB] = 8'hAF;
mem[16'h8ADC] = 8'h8A;
mem[16'h8ADD] = 8'h8D;
mem[16'h8ADE] = 8'hBC;
mem[16'h8ADF] = 8'h8A;
mem[16'h8AE0] = 8'h8C;
mem[16'h8AE1] = 8'h8F;
mem[16'h8AE2] = 8'h8A;
mem[16'h8AE3] = 8'h8C;
mem[16'h8AE4] = 8'h96;
mem[16'h8AE5] = 8'h8A;
mem[16'h8AE6] = 8'h8C;
mem[16'h8AE7] = 8'hA3;
mem[16'h8AE8] = 8'h8A;
mem[16'h8AE9] = 8'h8C;
mem[16'h8AEA] = 8'hB0;
mem[16'h8AEB] = 8'h8A;
mem[16'h8AEC] = 8'h8C;
mem[16'h8AED] = 8'hBD;
mem[16'h8AEE] = 8'h8A;
mem[16'h8AEF] = 8'h60;
mem[16'h8AF0] = 8'hA2;
mem[16'h8AF1] = 8'h00;
mem[16'h8AF2] = 8'hA4;
mem[16'h8AF3] = 8'h56;
mem[16'h8AF4] = 8'hB9;
mem[16'h8AF5] = 8'hD5;
mem[16'h8AF6] = 8'h8E;
mem[16'h8AF7] = 8'h85;
mem[16'h8AF8] = 8'h59;
mem[16'h8AF9] = 8'hB9;
mem[16'h8AFA] = 8'h95;
mem[16'h8AFB] = 8'h8F;
mem[16'h8AFC] = 8'h85;
mem[16'h8AFD] = 8'h5A;
mem[16'h8AFE] = 8'hA4;
mem[16'h8AFF] = 8'h57;
mem[16'h8B00] = 8'hB9;
mem[16'h8B01] = 8'h56;
mem[16'h8B02] = 8'h8D;
mem[16'h8B03] = 8'hA8;
mem[16'h8B04] = 8'hBD;
mem[16'h8B05] = 8'h38;
mem[16'h8B06] = 8'h81;
mem[16'h8B07] = 8'h29;
mem[16'h8B08] = 8'h80;
mem[16'h8B09] = 8'h85;
mem[16'h8B0A] = 8'h6D;
mem[16'h8B0B] = 8'hBD;
mem[16'h8B0C] = 8'h38;
mem[16'h8B0D] = 8'h81;
mem[16'h8B0E] = 8'h29;
mem[16'h8B0F] = 8'h7F;
mem[16'h8B10] = 8'h51;
mem[16'h8B11] = 8'h59;
mem[16'h8B12] = 8'h05;
mem[16'h8B13] = 8'h6D;
mem[16'h8B14] = 8'h91;
mem[16'h8B15] = 8'h59;
mem[16'h8B16] = 8'hE8;
mem[16'h8B17] = 8'hC8;
mem[16'h8B18] = 8'hBD;
mem[16'h8B19] = 8'h38;
mem[16'h8B1A] = 8'h81;
mem[16'h8B1B] = 8'h29;
mem[16'h8B1C] = 8'h7F;
mem[16'h8B1D] = 8'h51;
mem[16'h8B1E] = 8'h59;
mem[16'h8B1F] = 8'h05;
mem[16'h8B20] = 8'h6D;
mem[16'h8B21] = 8'h91;
mem[16'h8B22] = 8'h59;
mem[16'h8B23] = 8'hC8;
mem[16'h8B24] = 8'hE8;
mem[16'h8B25] = 8'hBD;
mem[16'h8B26] = 8'h38;
mem[16'h8B27] = 8'h81;
mem[16'h8B28] = 8'h29;
mem[16'h8B29] = 8'h7F;
mem[16'h8B2A] = 8'h51;
mem[16'h8B2B] = 8'h59;
mem[16'h8B2C] = 8'h05;
mem[16'h8B2D] = 8'h6D;
mem[16'h8B2E] = 8'h91;
mem[16'h8B2F] = 8'h59;
mem[16'h8B30] = 8'hE6;
mem[16'h8B31] = 8'h56;
mem[16'h8B32] = 8'hE8;
mem[16'h8B33] = 8'hE0;
mem[16'h8B34] = 8'h1B;
mem[16'h8B35] = 8'hB0;
mem[16'h8B36] = 8'h03;
mem[16'h8B37] = 8'h4C;
mem[16'h8B38] = 8'hF2;
mem[16'h8B39] = 8'h8A;
mem[16'h8B3A] = 8'h60;
mem[16'h8B3B] = 8'h8D;
mem[16'h8B3C] = 8'h05;
mem[16'h8B3D] = 8'h8B;
mem[16'h8B3E] = 8'h8D;
mem[16'h8B3F] = 8'h0C;
mem[16'h8B40] = 8'h8B;
mem[16'h8B41] = 8'h8D;
mem[16'h8B42] = 8'h19;
mem[16'h8B43] = 8'h8B;
mem[16'h8B44] = 8'h8D;
mem[16'h8B45] = 8'h26;
mem[16'h8B46] = 8'h8B;
mem[16'h8B47] = 8'h8C;
mem[16'h8B48] = 8'h06;
mem[16'h8B49] = 8'h8B;
mem[16'h8B4A] = 8'h8C;
mem[16'h8B4B] = 8'h0D;
mem[16'h8B4C] = 8'h8B;
mem[16'h8B4D] = 8'h8C;
mem[16'h8B4E] = 8'h1A;
mem[16'h8B4F] = 8'h8B;
mem[16'h8B50] = 8'h8C;
mem[16'h8B51] = 8'h27;
mem[16'h8B52] = 8'h8B;
mem[16'h8B53] = 8'h60;
mem[16'h8B54] = 8'hA2;
mem[16'h8B55] = 8'h00;
mem[16'h8B56] = 8'hA4;
mem[16'h8B57] = 8'h56;
mem[16'h8B58] = 8'hB9;
mem[16'h8B59] = 8'hD5;
mem[16'h8B5A] = 8'h8E;
mem[16'h8B5B] = 8'h85;
mem[16'h8B5C] = 8'h59;
mem[16'h8B5D] = 8'hB9;
mem[16'h8B5E] = 8'h95;
mem[16'h8B5F] = 8'h8F;
mem[16'h8B60] = 8'h85;
mem[16'h8B61] = 8'h5A;
mem[16'h8B62] = 8'hA0;
mem[16'h8B63] = 8'h26;
mem[16'h8B64] = 8'hBD;
mem[16'h8B65] = 8'hF3;
mem[16'h8B66] = 8'h4C;
mem[16'h8B67] = 8'h29;
mem[16'h8B68] = 8'h7F;
mem[16'h8B69] = 8'h51;
mem[16'h8B6A] = 8'h59;
mem[16'h8B6B] = 8'h91;
mem[16'h8B6C] = 8'h59;
mem[16'h8B6D] = 8'hE8;
mem[16'h8B6E] = 8'hC8;
mem[16'h8B6F] = 8'hBD;
mem[16'h8B70] = 8'hF3;
mem[16'h8B71] = 8'h4C;
mem[16'h8B72] = 8'h29;
mem[16'h8B73] = 8'h7F;
mem[16'h8B74] = 8'h51;
mem[16'h8B75] = 8'h59;
mem[16'h8B76] = 8'h91;
mem[16'h8B77] = 8'h59;
mem[16'h8B78] = 8'hE6;
mem[16'h8B79] = 8'h56;
mem[16'h8B7A] = 8'hE8;
mem[16'h8B7B] = 8'hE0;
mem[16'h8B7C] = 8'h1A;
mem[16'h8B7D] = 8'hB0;
mem[16'h8B7E] = 8'h03;
mem[16'h8B7F] = 8'h4C;
mem[16'h8B80] = 8'h56;
mem[16'h8B81] = 8'h8B;
mem[16'h8B82] = 8'h60;
mem[16'h8B83] = 8'hA9;
mem[16'h8B84] = 8'h92;
mem[16'h8B85] = 8'h85;
mem[16'h8B86] = 8'h59;
mem[16'h8B87] = 8'hA9;
mem[16'h8B88] = 8'h8B;
mem[16'h8B89] = 8'h85;
mem[16'h8B8A] = 8'h5A;
mem[16'h8B8B] = 8'h20;
mem[16'h8B8C] = 8'h8E;
mem[16'h8B8D] = 8'hFD;
mem[16'h8B8E] = 8'h20;
mem[16'h8B8F] = 8'hD5;
mem[16'h8B90] = 8'h67;
mem[16'h8B91] = 8'h60;
mem[16'h8B92] = 8'h84;
mem[16'h8B93] = 8'hC2;
mem[16'h8B94] = 8'hCC;
mem[16'h8B95] = 8'hCF;
mem[16'h8B96] = 8'hC1;
mem[16'h8B97] = 8'hC4;
mem[16'h8B98] = 8'hA0;
mem[16'h8B99] = 8'hD4;
mem[16'h8B9A] = 8'hC5;
mem[16'h8B9B] = 8'hD8;
mem[16'h8B9C] = 8'hD4;
mem[16'h8B9D] = 8'hAE;
mem[16'h8B9E] = 8'hB3;
mem[16'h8B9F] = 8'hB0;
mem[16'h8BA0] = 8'hB0;
mem[16'h8BA1] = 8'hAC;
mem[16'h8BA2] = 8'hC1;
mem[16'h8BA3] = 8'hA4;
mem[16'h8BA4] = 8'hB3;
mem[16'h8BA5] = 8'hB0;
mem[16'h8BA6] = 8'hB0;
mem[16'h8BA7] = 8'h00;
mem[16'h8BA8] = 8'hA2;
mem[16'h8BA9] = 8'h00;
mem[16'h8BAA] = 8'hA4;
mem[16'h8BAB] = 8'h56;
mem[16'h8BAC] = 8'hB9;
mem[16'h8BAD] = 8'hD5;
mem[16'h8BAE] = 8'h8E;
mem[16'h8BAF] = 8'h85;
mem[16'h8BB0] = 8'h59;
mem[16'h8BB1] = 8'hB9;
mem[16'h8BB2] = 8'h95;
mem[16'h8BB3] = 8'h8F;
mem[16'h8BB4] = 8'h85;
mem[16'h8BB5] = 8'h5A;
mem[16'h8BB6] = 8'hA4;
mem[16'h8BB7] = 8'h57;
mem[16'h8BB8] = 8'hB9;
mem[16'h8BB9] = 8'h3E;
mem[16'h8BBA] = 8'h8C;
mem[16'h8BBB] = 8'h85;
mem[16'h8BBC] = 8'h5C;
mem[16'h8BBD] = 8'hB9;
mem[16'h8BBE] = 8'h56;
mem[16'h8BBF] = 8'h8D;
mem[16'h8BC0] = 8'hA8;
mem[16'h8BC1] = 8'hBD;
mem[16'h8BC2] = 8'h08;
mem[16'h8BC3] = 8'h5F;
mem[16'h8BC4] = 8'h29;
mem[16'h8BC5] = 8'h80;
mem[16'h8BC6] = 8'h85;
mem[16'h8BC7] = 8'h6D;
mem[16'h8BC8] = 8'hBD;
mem[16'h8BC9] = 8'h08;
mem[16'h8BCA] = 8'h5F;
mem[16'h8BCB] = 8'h29;
mem[16'h8BCC] = 8'h7F;
mem[16'h8BCD] = 8'h85;
mem[16'h8BCE] = 8'h66;
mem[16'h8BCF] = 8'hE8;
mem[16'h8BD0] = 8'hBD;
mem[16'h8BD1] = 8'h08;
mem[16'h8BD2] = 8'h5F;
mem[16'h8BD3] = 8'h29;
mem[16'h8BD4] = 8'h7F;
mem[16'h8BD5] = 8'h85;
mem[16'h8BD6] = 8'h67;
mem[16'h8BD7] = 8'hA9;
mem[16'h8BD8] = 8'h00;
mem[16'h8BD9] = 8'h85;
mem[16'h8BDA] = 8'h68;
mem[16'h8BDB] = 8'h85;
mem[16'h8BDC] = 8'h6A;
mem[16'h8BDD] = 8'hA5;
mem[16'h8BDE] = 8'h5C;
mem[16'h8BDF] = 8'hC9;
mem[16'h8BE0] = 8'h01;
mem[16'h8BE1] = 8'hF0;
mem[16'h8BE2] = 8'h23;
mem[16'h8BE3] = 8'h46;
mem[16'h8BE4] = 8'h67;
mem[16'h8BE5] = 8'h66;
mem[16'h8BE6] = 8'h6A;
mem[16'h8BE7] = 8'h46;
mem[16'h8BE8] = 8'h66;
mem[16'h8BE9] = 8'h66;
mem[16'h8BEA] = 8'h68;
mem[16'h8BEB] = 8'h06;
mem[16'h8BEC] = 8'h5C;
mem[16'h8BED] = 8'h24;
mem[16'h8BEE] = 8'h5C;
mem[16'h8BEF] = 8'h10;
mem[16'h8BF0] = 8'hF2;
mem[16'h8BF1] = 8'h46;
mem[16'h8BF2] = 8'h68;
mem[16'h8BF3] = 8'hA5;
mem[16'h8BF4] = 8'h6A;
mem[16'h8BF5] = 8'h4A;
mem[16'h8BF6] = 8'h05;
mem[16'h8BF7] = 8'h66;
mem[16'h8BF8] = 8'h85;
mem[16'h8BF9] = 8'h6A;
mem[16'h8BFA] = 8'hA5;
mem[16'h8BFB] = 8'h68;
mem[16'h8BFC] = 8'h85;
mem[16'h8BFD] = 8'h66;
mem[16'h8BFE] = 8'hA5;
mem[16'h8BFF] = 8'h67;
mem[16'h8C00] = 8'h85;
mem[16'h8C01] = 8'h68;
mem[16'h8C02] = 8'hA5;
mem[16'h8C03] = 8'h6A;
mem[16'h8C04] = 8'h85;
mem[16'h8C05] = 8'h67;
mem[16'h8C06] = 8'hA5;
mem[16'h8C07] = 8'h66;
mem[16'h8C08] = 8'h05;
mem[16'h8C09] = 8'h6D;
mem[16'h8C0A] = 8'h51;
mem[16'h8C0B] = 8'h59;
mem[16'h8C0C] = 8'h91;
mem[16'h8C0D] = 8'h59;
mem[16'h8C0E] = 8'hC8;
mem[16'h8C0F] = 8'hA5;
mem[16'h8C10] = 8'h67;
mem[16'h8C11] = 8'h05;
mem[16'h8C12] = 8'h6D;
mem[16'h8C13] = 8'h51;
mem[16'h8C14] = 8'h59;
mem[16'h8C15] = 8'h91;
mem[16'h8C16] = 8'h59;
mem[16'h8C17] = 8'hC8;
mem[16'h8C18] = 8'hA5;
mem[16'h8C19] = 8'h68;
mem[16'h8C1A] = 8'h05;
mem[16'h8C1B] = 8'h6D;
mem[16'h8C1C] = 8'h51;
mem[16'h8C1D] = 8'h59;
mem[16'h8C1E] = 8'h91;
mem[16'h8C1F] = 8'h59;
mem[16'h8C20] = 8'hE6;
mem[16'h8C21] = 8'h56;
mem[16'h8C22] = 8'hE8;
mem[16'h8C23] = 8'hE0;
mem[16'h8C24] = 8'h16;
mem[16'h8C25] = 8'hB0;
mem[16'h8C26] = 8'h03;
mem[16'h8C27] = 8'h4C;
mem[16'h8C28] = 8'hAA;
mem[16'h8C29] = 8'h8B;
mem[16'h8C2A] = 8'h60;
mem[16'h8C2B] = 8'h8D;
mem[16'h8C2C] = 8'hC2;
mem[16'h8C2D] = 8'h8B;
mem[16'h8C2E] = 8'h8D;
mem[16'h8C2F] = 8'hC9;
mem[16'h8C30] = 8'h8B;
mem[16'h8C31] = 8'h8D;
mem[16'h8C32] = 8'hD1;
mem[16'h8C33] = 8'h8B;
mem[16'h8C34] = 8'h8C;
mem[16'h8C35] = 8'hC3;
mem[16'h8C36] = 8'h8B;
mem[16'h8C37] = 8'h8C;
mem[16'h8C38] = 8'hCA;
mem[16'h8C39] = 8'h8B;
mem[16'h8C3A] = 8'h8C;
mem[16'h8C3B] = 8'hD2;
mem[16'h8C3C] = 8'h8B;
mem[16'h8C3D] = 8'h60;
mem[16'h8C3E] = 8'h01;
mem[16'h8C3F] = 8'h02;
mem[16'h8C40] = 8'h04;
mem[16'h8C41] = 8'h08;
mem[16'h8C42] = 8'h10;
mem[16'h8C43] = 8'h20;
mem[16'h8C44] = 8'h40;
mem[16'h8C45] = 8'h01;
mem[16'h8C46] = 8'h02;
mem[16'h8C47] = 8'h04;
mem[16'h8C48] = 8'h08;
mem[16'h8C49] = 8'h10;
mem[16'h8C4A] = 8'h20;
mem[16'h8C4B] = 8'h40;
mem[16'h8C4C] = 8'h01;
mem[16'h8C4D] = 8'h02;
mem[16'h8C4E] = 8'h04;
mem[16'h8C4F] = 8'h08;
mem[16'h8C50] = 8'h10;
mem[16'h8C51] = 8'h20;
mem[16'h8C52] = 8'h40;
mem[16'h8C53] = 8'h01;
mem[16'h8C54] = 8'h02;
mem[16'h8C55] = 8'h04;
mem[16'h8C56] = 8'h08;
mem[16'h8C57] = 8'h10;
mem[16'h8C58] = 8'h20;
mem[16'h8C59] = 8'h40;
mem[16'h8C5A] = 8'h01;
mem[16'h8C5B] = 8'h02;
mem[16'h8C5C] = 8'h04;
mem[16'h8C5D] = 8'h08;
mem[16'h8C5E] = 8'h10;
mem[16'h8C5F] = 8'h20;
mem[16'h8C60] = 8'h40;
mem[16'h8C61] = 8'h01;
mem[16'h8C62] = 8'h02;
mem[16'h8C63] = 8'h04;
mem[16'h8C64] = 8'h08;
mem[16'h8C65] = 8'h10;
mem[16'h8C66] = 8'h20;
mem[16'h8C67] = 8'h40;
mem[16'h8C68] = 8'h01;
mem[16'h8C69] = 8'h02;
mem[16'h8C6A] = 8'h04;
mem[16'h8C6B] = 8'h08;
mem[16'h8C6C] = 8'h10;
mem[16'h8C6D] = 8'h20;
mem[16'h8C6E] = 8'h40;
mem[16'h8C6F] = 8'h01;
mem[16'h8C70] = 8'h02;
mem[16'h8C71] = 8'h04;
mem[16'h8C72] = 8'h08;
mem[16'h8C73] = 8'h10;
mem[16'h8C74] = 8'h20;
mem[16'h8C75] = 8'h40;
mem[16'h8C76] = 8'h01;
mem[16'h8C77] = 8'h02;
mem[16'h8C78] = 8'h04;
mem[16'h8C79] = 8'h08;
mem[16'h8C7A] = 8'h10;
mem[16'h8C7B] = 8'h20;
mem[16'h8C7C] = 8'h40;
mem[16'h8C7D] = 8'h01;
mem[16'h8C7E] = 8'h02;
mem[16'h8C7F] = 8'h04;
mem[16'h8C80] = 8'h08;
mem[16'h8C81] = 8'h10;
mem[16'h8C82] = 8'h20;
mem[16'h8C83] = 8'h40;
mem[16'h8C84] = 8'h01;
mem[16'h8C85] = 8'h02;
mem[16'h8C86] = 8'h04;
mem[16'h8C87] = 8'h08;
mem[16'h8C88] = 8'h10;
mem[16'h8C89] = 8'h20;
mem[16'h8C8A] = 8'h40;
mem[16'h8C8B] = 8'h01;
mem[16'h8C8C] = 8'h02;
mem[16'h8C8D] = 8'h04;
mem[16'h8C8E] = 8'h08;
mem[16'h8C8F] = 8'h10;
mem[16'h8C90] = 8'h20;
mem[16'h8C91] = 8'h40;
mem[16'h8C92] = 8'h01;
mem[16'h8C93] = 8'h02;
mem[16'h8C94] = 8'h04;
mem[16'h8C95] = 8'h08;
mem[16'h8C96] = 8'h10;
mem[16'h8C97] = 8'h20;
mem[16'h8C98] = 8'h40;
mem[16'h8C99] = 8'h01;
mem[16'h8C9A] = 8'h02;
mem[16'h8C9B] = 8'h04;
mem[16'h8C9C] = 8'h08;
mem[16'h8C9D] = 8'h10;
mem[16'h8C9E] = 8'h20;
mem[16'h8C9F] = 8'h40;
mem[16'h8CA0] = 8'h01;
mem[16'h8CA1] = 8'h02;
mem[16'h8CA2] = 8'h04;
mem[16'h8CA3] = 8'h08;
mem[16'h8CA4] = 8'h10;
mem[16'h8CA5] = 8'h20;
mem[16'h8CA6] = 8'h40;
mem[16'h8CA7] = 8'h01;
mem[16'h8CA8] = 8'h02;
mem[16'h8CA9] = 8'h04;
mem[16'h8CAA] = 8'h08;
mem[16'h8CAB] = 8'h10;
mem[16'h8CAC] = 8'h20;
mem[16'h8CAD] = 8'h40;
mem[16'h8CAE] = 8'h01;
mem[16'h8CAF] = 8'h02;
mem[16'h8CB0] = 8'h04;
mem[16'h8CB1] = 8'h08;
mem[16'h8CB2] = 8'h10;
mem[16'h8CB3] = 8'h20;
mem[16'h8CB4] = 8'h40;
mem[16'h8CB5] = 8'h01;
mem[16'h8CB6] = 8'h02;
mem[16'h8CB7] = 8'h04;
mem[16'h8CB8] = 8'h08;
mem[16'h8CB9] = 8'h10;
mem[16'h8CBA] = 8'h20;
mem[16'h8CBB] = 8'h40;
mem[16'h8CBC] = 8'h01;
mem[16'h8CBD] = 8'h02;
mem[16'h8CBE] = 8'h04;
mem[16'h8CBF] = 8'h08;
mem[16'h8CC0] = 8'h10;
mem[16'h8CC1] = 8'h20;
mem[16'h8CC2] = 8'h40;
mem[16'h8CC3] = 8'h01;
mem[16'h8CC4] = 8'h02;
mem[16'h8CC5] = 8'h04;
mem[16'h8CC6] = 8'h08;
mem[16'h8CC7] = 8'h10;
mem[16'h8CC8] = 8'h20;
mem[16'h8CC9] = 8'h40;
mem[16'h8CCA] = 8'h01;
mem[16'h8CCB] = 8'h02;
mem[16'h8CCC] = 8'h04;
mem[16'h8CCD] = 8'h08;
mem[16'h8CCE] = 8'h10;
mem[16'h8CCF] = 8'h20;
mem[16'h8CD0] = 8'h40;
mem[16'h8CD1] = 8'h01;
mem[16'h8CD2] = 8'h02;
mem[16'h8CD3] = 8'h04;
mem[16'h8CD4] = 8'h08;
mem[16'h8CD5] = 8'h10;
mem[16'h8CD6] = 8'h20;
mem[16'h8CD7] = 8'h40;
mem[16'h8CD8] = 8'h01;
mem[16'h8CD9] = 8'h02;
mem[16'h8CDA] = 8'h04;
mem[16'h8CDB] = 8'h08;
mem[16'h8CDC] = 8'h10;
mem[16'h8CDD] = 8'h20;
mem[16'h8CDE] = 8'h40;
mem[16'h8CDF] = 8'h01;
mem[16'h8CE0] = 8'h02;
mem[16'h8CE1] = 8'h04;
mem[16'h8CE2] = 8'h08;
mem[16'h8CE3] = 8'h10;
mem[16'h8CE4] = 8'h20;
mem[16'h8CE5] = 8'h40;
mem[16'h8CE6] = 8'h01;
mem[16'h8CE7] = 8'h02;
mem[16'h8CE8] = 8'h04;
mem[16'h8CE9] = 8'h08;
mem[16'h8CEA] = 8'h10;
mem[16'h8CEB] = 8'h20;
mem[16'h8CEC] = 8'h40;
mem[16'h8CED] = 8'h01;
mem[16'h8CEE] = 8'h02;
mem[16'h8CEF] = 8'h04;
mem[16'h8CF0] = 8'h08;
mem[16'h8CF1] = 8'h10;
mem[16'h8CF2] = 8'h20;
mem[16'h8CF3] = 8'h40;
mem[16'h8CF4] = 8'h01;
mem[16'h8CF5] = 8'h02;
mem[16'h8CF6] = 8'h04;
mem[16'h8CF7] = 8'h08;
mem[16'h8CF8] = 8'h10;
mem[16'h8CF9] = 8'h20;
mem[16'h8CFA] = 8'h40;
mem[16'h8CFB] = 8'h01;
mem[16'h8CFC] = 8'h02;
mem[16'h8CFD] = 8'h04;
mem[16'h8CFE] = 8'h08;
mem[16'h8CFF] = 8'h10;
mem[16'h8D00] = 8'h20;
mem[16'h8D01] = 8'h40;
mem[16'h8D02] = 8'h01;
mem[16'h8D03] = 8'h02;
mem[16'h8D04] = 8'h04;
mem[16'h8D05] = 8'h08;
mem[16'h8D06] = 8'h10;
mem[16'h8D07] = 8'h20;
mem[16'h8D08] = 8'h40;
mem[16'h8D09] = 8'h01;
mem[16'h8D0A] = 8'h02;
mem[16'h8D0B] = 8'h04;
mem[16'h8D0C] = 8'h08;
mem[16'h8D0D] = 8'h10;
mem[16'h8D0E] = 8'h20;
mem[16'h8D0F] = 8'h40;
mem[16'h8D10] = 8'h01;
mem[16'h8D11] = 8'h02;
mem[16'h8D12] = 8'h04;
mem[16'h8D13] = 8'h08;
mem[16'h8D14] = 8'h10;
mem[16'h8D15] = 8'h20;
mem[16'h8D16] = 8'h40;
mem[16'h8D17] = 8'h01;
mem[16'h8D18] = 8'h02;
mem[16'h8D19] = 8'h04;
mem[16'h8D1A] = 8'h08;
mem[16'h8D1B] = 8'h10;
mem[16'h8D1C] = 8'h20;
mem[16'h8D1D] = 8'h40;
mem[16'h8D1E] = 8'h01;
mem[16'h8D1F] = 8'h02;
mem[16'h8D20] = 8'h04;
mem[16'h8D21] = 8'h08;
mem[16'h8D22] = 8'h10;
mem[16'h8D23] = 8'h20;
mem[16'h8D24] = 8'h40;
mem[16'h8D25] = 8'h01;
mem[16'h8D26] = 8'h02;
mem[16'h8D27] = 8'h04;
mem[16'h8D28] = 8'h08;
mem[16'h8D29] = 8'h10;
mem[16'h8D2A] = 8'h20;
mem[16'h8D2B] = 8'h40;
mem[16'h8D2C] = 8'h01;
mem[16'h8D2D] = 8'h02;
mem[16'h8D2E] = 8'h04;
mem[16'h8D2F] = 8'h08;
mem[16'h8D30] = 8'h10;
mem[16'h8D31] = 8'h20;
mem[16'h8D32] = 8'h40;
mem[16'h8D33] = 8'h01;
mem[16'h8D34] = 8'h02;
mem[16'h8D35] = 8'h04;
mem[16'h8D36] = 8'h08;
mem[16'h8D37] = 8'h10;
mem[16'h8D38] = 8'h20;
mem[16'h8D39] = 8'h40;
mem[16'h8D3A] = 8'h01;
mem[16'h8D3B] = 8'h02;
mem[16'h8D3C] = 8'h04;
mem[16'h8D3D] = 8'h08;
mem[16'h8D3E] = 8'h10;
mem[16'h8D3F] = 8'h20;
mem[16'h8D40] = 8'h40;
mem[16'h8D41] = 8'h01;
mem[16'h8D42] = 8'h02;
mem[16'h8D43] = 8'h04;
mem[16'h8D44] = 8'h08;
mem[16'h8D45] = 8'h10;
mem[16'h8D46] = 8'h20;
mem[16'h8D47] = 8'h40;
mem[16'h8D48] = 8'h01;
mem[16'h8D49] = 8'h02;
mem[16'h8D4A] = 8'h04;
mem[16'h8D4B] = 8'h08;
mem[16'h8D4C] = 8'h10;
mem[16'h8D4D] = 8'h20;
mem[16'h8D4E] = 8'h40;
mem[16'h8D4F] = 8'h01;
mem[16'h8D50] = 8'h02;
mem[16'h8D51] = 8'h04;
mem[16'h8D52] = 8'h08;
mem[16'h8D53] = 8'h10;
mem[16'h8D54] = 8'h20;
mem[16'h8D55] = 8'h40;
mem[16'h8D56] = 8'h00;
mem[16'h8D57] = 8'h00;
mem[16'h8D58] = 8'h00;
mem[16'h8D59] = 8'h00;
mem[16'h8D5A] = 8'h00;
mem[16'h8D5B] = 8'h00;
mem[16'h8D5C] = 8'h00;
mem[16'h8D5D] = 8'h01;
mem[16'h8D5E] = 8'h01;
mem[16'h8D5F] = 8'h01;
mem[16'h8D60] = 8'h01;
mem[16'h8D61] = 8'h01;
mem[16'h8D62] = 8'h01;
mem[16'h8D63] = 8'h01;
mem[16'h8D64] = 8'h02;
mem[16'h8D65] = 8'h02;
mem[16'h8D66] = 8'h02;
mem[16'h8D67] = 8'h02;
mem[16'h8D68] = 8'h02;
mem[16'h8D69] = 8'h02;
mem[16'h8D6A] = 8'h02;
mem[16'h8D6B] = 8'h03;
mem[16'h8D6C] = 8'h03;
mem[16'h8D6D] = 8'h03;
mem[16'h8D6E] = 8'h03;
mem[16'h8D6F] = 8'h03;
mem[16'h8D70] = 8'h03;
mem[16'h8D71] = 8'h03;
mem[16'h8D72] = 8'h04;
mem[16'h8D73] = 8'h04;
mem[16'h8D74] = 8'h04;
mem[16'h8D75] = 8'h04;
mem[16'h8D76] = 8'h04;
mem[16'h8D77] = 8'h04;
mem[16'h8D78] = 8'h04;
mem[16'h8D79] = 8'h05;
mem[16'h8D7A] = 8'h05;
mem[16'h8D7B] = 8'h05;
mem[16'h8D7C] = 8'h05;
mem[16'h8D7D] = 8'h05;
mem[16'h8D7E] = 8'h05;
mem[16'h8D7F] = 8'h05;
mem[16'h8D80] = 8'h06;
mem[16'h8D81] = 8'h06;
mem[16'h8D82] = 8'h06;
mem[16'h8D83] = 8'h06;
mem[16'h8D84] = 8'h06;
mem[16'h8D85] = 8'h06;
mem[16'h8D86] = 8'h06;
mem[16'h8D87] = 8'h07;
mem[16'h8D88] = 8'h07;
mem[16'h8D89] = 8'h07;
mem[16'h8D8A] = 8'h07;
mem[16'h8D8B] = 8'h07;
mem[16'h8D8C] = 8'h07;
mem[16'h8D8D] = 8'h07;
mem[16'h8D8E] = 8'h08;
mem[16'h8D8F] = 8'h08;
mem[16'h8D90] = 8'h08;
mem[16'h8D91] = 8'h08;
mem[16'h8D92] = 8'h08;
mem[16'h8D93] = 8'h08;
mem[16'h8D94] = 8'h08;
mem[16'h8D95] = 8'h09;
mem[16'h8D96] = 8'h09;
mem[16'h8D97] = 8'h09;
mem[16'h8D98] = 8'h09;
mem[16'h8D99] = 8'h09;
mem[16'h8D9A] = 8'h09;
mem[16'h8D9B] = 8'h09;
mem[16'h8D9C] = 8'h0A;
mem[16'h8D9D] = 8'h0A;
mem[16'h8D9E] = 8'h0A;
mem[16'h8D9F] = 8'h0A;
mem[16'h8DA0] = 8'h0A;
mem[16'h8DA1] = 8'h0A;
mem[16'h8DA2] = 8'h0A;
mem[16'h8DA3] = 8'h0B;
mem[16'h8DA4] = 8'h0B;
mem[16'h8DA5] = 8'h0B;
mem[16'h8DA6] = 8'h0B;
mem[16'h8DA7] = 8'h0B;
mem[16'h8DA8] = 8'h0B;
mem[16'h8DA9] = 8'h0B;
mem[16'h8DAA] = 8'h0C;
mem[16'h8DAB] = 8'h0C;
mem[16'h8DAC] = 8'h0C;
mem[16'h8DAD] = 8'h0C;
mem[16'h8DAE] = 8'h0C;
mem[16'h8DAF] = 8'h0C;
mem[16'h8DB0] = 8'h0C;
mem[16'h8DB1] = 8'h0D;
mem[16'h8DB2] = 8'h0D;
mem[16'h8DB3] = 8'h0D;
mem[16'h8DB4] = 8'h0D;
mem[16'h8DB5] = 8'h0D;
mem[16'h8DB6] = 8'h0D;
mem[16'h8DB7] = 8'h0D;
mem[16'h8DB8] = 8'h0E;
mem[16'h8DB9] = 8'h0E;
mem[16'h8DBA] = 8'h0E;
mem[16'h8DBB] = 8'h0E;
mem[16'h8DBC] = 8'h0E;
mem[16'h8DBD] = 8'h0E;
mem[16'h8DBE] = 8'h0E;
mem[16'h8DBF] = 8'h0F;
mem[16'h8DC0] = 8'h0F;
mem[16'h8DC1] = 8'h0F;
mem[16'h8DC2] = 8'h0F;
mem[16'h8DC3] = 8'h0F;
mem[16'h8DC4] = 8'h0F;
mem[16'h8DC5] = 8'h0F;
mem[16'h8DC6] = 8'h10;
mem[16'h8DC7] = 8'h10;
mem[16'h8DC8] = 8'h10;
mem[16'h8DC9] = 8'h10;
mem[16'h8DCA] = 8'h10;
mem[16'h8DCB] = 8'h10;
mem[16'h8DCC] = 8'h10;
mem[16'h8DCD] = 8'h11;
mem[16'h8DCE] = 8'h11;
mem[16'h8DCF] = 8'h11;
mem[16'h8DD0] = 8'h11;
mem[16'h8DD1] = 8'h11;
mem[16'h8DD2] = 8'h11;
mem[16'h8DD3] = 8'h11;
mem[16'h8DD4] = 8'h12;
mem[16'h8DD5] = 8'h12;
mem[16'h8DD6] = 8'h12;
mem[16'h8DD7] = 8'h12;
mem[16'h8DD8] = 8'h12;
mem[16'h8DD9] = 8'h12;
mem[16'h8DDA] = 8'h12;
mem[16'h8DDB] = 8'h13;
mem[16'h8DDC] = 8'h13;
mem[16'h8DDD] = 8'h13;
mem[16'h8DDE] = 8'h13;
mem[16'h8DDF] = 8'h13;
mem[16'h8DE0] = 8'h13;
mem[16'h8DE1] = 8'h13;
mem[16'h8DE2] = 8'h14;
mem[16'h8DE3] = 8'h14;
mem[16'h8DE4] = 8'h14;
mem[16'h8DE5] = 8'h14;
mem[16'h8DE6] = 8'h14;
mem[16'h8DE7] = 8'h14;
mem[16'h8DE8] = 8'h14;
mem[16'h8DE9] = 8'h15;
mem[16'h8DEA] = 8'h15;
mem[16'h8DEB] = 8'h15;
mem[16'h8DEC] = 8'h15;
mem[16'h8DED] = 8'h15;
mem[16'h8DEE] = 8'h15;
mem[16'h8DEF] = 8'h15;
mem[16'h8DF0] = 8'h16;
mem[16'h8DF1] = 8'h16;
mem[16'h8DF2] = 8'h16;
mem[16'h8DF3] = 8'h16;
mem[16'h8DF4] = 8'h16;
mem[16'h8DF5] = 8'h16;
mem[16'h8DF6] = 8'h16;
mem[16'h8DF7] = 8'h17;
mem[16'h8DF8] = 8'h17;
mem[16'h8DF9] = 8'h17;
mem[16'h8DFA] = 8'h17;
mem[16'h8DFB] = 8'h17;
mem[16'h8DFC] = 8'h17;
mem[16'h8DFD] = 8'h17;
mem[16'h8DFE] = 8'h18;
mem[16'h8DFF] = 8'h18;
mem[16'h8E00] = 8'h18;
mem[16'h8E01] = 8'h18;
mem[16'h8E02] = 8'h18;
mem[16'h8E03] = 8'h18;
mem[16'h8E04] = 8'h18;
mem[16'h8E05] = 8'h19;
mem[16'h8E06] = 8'h19;
mem[16'h8E07] = 8'h19;
mem[16'h8E08] = 8'h19;
mem[16'h8E09] = 8'h19;
mem[16'h8E0A] = 8'h19;
mem[16'h8E0B] = 8'h19;
mem[16'h8E0C] = 8'h1A;
mem[16'h8E0D] = 8'h1A;
mem[16'h8E0E] = 8'h1A;
mem[16'h8E0F] = 8'h1A;
mem[16'h8E10] = 8'h1A;
mem[16'h8E11] = 8'h1A;
mem[16'h8E12] = 8'h1A;
mem[16'h8E13] = 8'h1B;
mem[16'h8E14] = 8'h1B;
mem[16'h8E15] = 8'h1B;
mem[16'h8E16] = 8'h1B;
mem[16'h8E17] = 8'h1B;
mem[16'h8E18] = 8'h1B;
mem[16'h8E19] = 8'h1B;
mem[16'h8E1A] = 8'h1C;
mem[16'h8E1B] = 8'h1C;
mem[16'h8E1C] = 8'h1C;
mem[16'h8E1D] = 8'h1C;
mem[16'h8E1E] = 8'h1C;
mem[16'h8E1F] = 8'h1C;
mem[16'h8E20] = 8'h1C;
mem[16'h8E21] = 8'h1D;
mem[16'h8E22] = 8'h1D;
mem[16'h8E23] = 8'h1D;
mem[16'h8E24] = 8'h1D;
mem[16'h8E25] = 8'h1D;
mem[16'h8E26] = 8'h1D;
mem[16'h8E27] = 8'h1D;
mem[16'h8E28] = 8'h1E;
mem[16'h8E29] = 8'h1E;
mem[16'h8E2A] = 8'h1E;
mem[16'h8E2B] = 8'h1E;
mem[16'h8E2C] = 8'h1E;
mem[16'h8E2D] = 8'h1E;
mem[16'h8E2E] = 8'h1E;
mem[16'h8E2F] = 8'h1F;
mem[16'h8E30] = 8'h1F;
mem[16'h8E31] = 8'h1F;
mem[16'h8E32] = 8'h1F;
mem[16'h8E33] = 8'h1F;
mem[16'h8E34] = 8'h1F;
mem[16'h8E35] = 8'h1F;
mem[16'h8E36] = 8'h20;
mem[16'h8E37] = 8'h20;
mem[16'h8E38] = 8'h20;
mem[16'h8E39] = 8'h20;
mem[16'h8E3A] = 8'h20;
mem[16'h8E3B] = 8'h20;
mem[16'h8E3C] = 8'h20;
mem[16'h8E3D] = 8'h21;
mem[16'h8E3E] = 8'h21;
mem[16'h8E3F] = 8'h21;
mem[16'h8E40] = 8'h21;
mem[16'h8E41] = 8'h21;
mem[16'h8E42] = 8'h21;
mem[16'h8E43] = 8'h21;
mem[16'h8E44] = 8'h22;
mem[16'h8E45] = 8'h22;
mem[16'h8E46] = 8'h22;
mem[16'h8E47] = 8'h22;
mem[16'h8E48] = 8'h22;
mem[16'h8E49] = 8'h22;
mem[16'h8E4A] = 8'h22;
mem[16'h8E4B] = 8'h23;
mem[16'h8E4C] = 8'h23;
mem[16'h8E4D] = 8'h23;
mem[16'h8E4E] = 8'h23;
mem[16'h8E4F] = 8'h23;
mem[16'h8E50] = 8'h23;
mem[16'h8E51] = 8'h23;
mem[16'h8E52] = 8'h24;
mem[16'h8E53] = 8'h24;
mem[16'h8E54] = 8'h24;
mem[16'h8E55] = 8'h24;
mem[16'h8E56] = 8'h24;
mem[16'h8E57] = 8'h24;
mem[16'h8E58] = 8'h24;
mem[16'h8E59] = 8'h25;
mem[16'h8E5A] = 8'h25;
mem[16'h8E5B] = 8'h25;
mem[16'h8E5C] = 8'h25;
mem[16'h8E5D] = 8'h25;
mem[16'h8E5E] = 8'h25;
mem[16'h8E5F] = 8'h25;
mem[16'h8E60] = 8'h26;
mem[16'h8E61] = 8'h26;
mem[16'h8E62] = 8'h26;
mem[16'h8E63] = 8'h26;
mem[16'h8E64] = 8'h26;
mem[16'h8E65] = 8'h26;
mem[16'h8E66] = 8'h26;
mem[16'h8E67] = 8'h27;
mem[16'h8E68] = 8'h27;
mem[16'h8E69] = 8'h27;
mem[16'h8E6A] = 8'h27;
mem[16'h8E6B] = 8'h27;
mem[16'h8E6C] = 8'h27;
mem[16'h8E6D] = 8'h27;
mem[16'h8E6E] = 8'h24;
mem[16'h8E6F] = 8'h24;
mem[16'h8E70] = 8'h24;
mem[16'h8E71] = 8'h25;
mem[16'h8E72] = 8'h25;
mem[16'h8E73] = 8'h25;
mem[16'h8E74] = 8'h25;
mem[16'h8E75] = 8'h25;
mem[16'h8E76] = 8'h25;
mem[16'h8E77] = 8'h25;
mem[16'h8E78] = 8'h26;
mem[16'h8E79] = 8'h26;
mem[16'h8E7A] = 8'h26;
mem[16'h8E7B] = 8'h26;
mem[16'h8E7C] = 8'h26;
mem[16'h8E7D] = 8'h26;
mem[16'h8E7E] = 8'h26;
mem[16'h8E7F] = 8'h27;
mem[16'h8E80] = 8'h27;
mem[16'h8E81] = 8'h27;
mem[16'h8E82] = 8'h27;
mem[16'h8E83] = 8'h27;
mem[16'h8E84] = 8'h27;
mem[16'h8E85] = 8'h27;
mem[16'h8E86] = 8'h28;
mem[16'h8E87] = 8'h28;
mem[16'h8E88] = 8'h28;
mem[16'h8E89] = 8'h28;
mem[16'h8E8A] = 8'h28;
mem[16'h8E8B] = 8'h28;
mem[16'h8E8C] = 8'h28;
mem[16'h8E8D] = 8'h29;
mem[16'h8E8E] = 8'h29;
mem[16'h8E8F] = 8'h29;
mem[16'h8E90] = 8'h29;
mem[16'h8E91] = 8'h29;
mem[16'h8E92] = 8'h29;
mem[16'h8E93] = 8'h29;
mem[16'h8E94] = 8'h00;
mem[16'h8E95] = 8'h00;
mem[16'h8E96] = 8'h01;
mem[16'h8E97] = 8'h00;
mem[16'h8E98] = 8'h02;
mem[16'h8E99] = 8'h00;
mem[16'h8E9A] = 8'h00;
mem[16'h8E9B] = 8'h00;
mem[16'h8E9C] = 8'h03;
mem[16'h8E9D] = 8'h00;
mem[16'h8E9E] = 8'h00;
mem[16'h8E9F] = 8'h00;
mem[16'h8EA0] = 8'h00;
mem[16'h8EA1] = 8'h00;
mem[16'h8EA2] = 8'h00;
mem[16'h8EA3] = 8'h00;
mem[16'h8EA4] = 8'h04;
mem[16'h8EA5] = 8'h00;
mem[16'h8EA6] = 8'h00;
mem[16'h8EA7] = 8'h00;
mem[16'h8EA8] = 8'h00;
mem[16'h8EA9] = 8'h00;
mem[16'h8EAA] = 8'h00;
mem[16'h8EAB] = 8'h00;
mem[16'h8EAC] = 8'h00;
mem[16'h8EAD] = 8'h00;
mem[16'h8EAE] = 8'h00;
mem[16'h8EAF] = 8'h00;
mem[16'h8EB0] = 8'h00;
mem[16'h8EB1] = 8'h00;
mem[16'h8EB2] = 8'h00;
mem[16'h8EB3] = 8'h00;
mem[16'h8EB4] = 8'h05;
mem[16'h8EB5] = 8'h00;
mem[16'h8EB6] = 8'hA2;
mem[16'h8EB7] = 8'hE6;
mem[16'h8EB8] = 8'h9A;
mem[16'h8EB9] = 8'hA9;
mem[16'h8EBA] = 8'h00;
mem[16'h8EBB] = 8'hA2;
mem[16'h8EBC] = 8'h16;
mem[16'h8EBD] = 8'hA0;
mem[16'h8EBE] = 8'h00;
mem[16'h8EBF] = 8'h78;
mem[16'h8EC0] = 8'h4C;
mem[16'h8EC1] = 8'h0B;
mem[16'h8EC2] = 8'h65;
mem[16'h8EC3] = 8'h00;
mem[16'h8EC4] = 8'h00;
mem[16'h8EC5] = 8'h00;
mem[16'h8EC6] = 8'h00;
mem[16'h8EC7] = 8'h00;
mem[16'h8EC8] = 8'h00;
mem[16'h8EC9] = 8'h00;
mem[16'h8ECA] = 8'h00;
mem[16'h8ECB] = 8'h00;
mem[16'h8ECC] = 8'h00;
mem[16'h8ECD] = 8'h00;
mem[16'h8ECE] = 8'h00;
mem[16'h8ECF] = 8'h00;
mem[16'h8ED0] = 8'h00;
mem[16'h8ED1] = 8'h00;
mem[16'h8ED2] = 8'h00;
mem[16'h8ED3] = 8'h00;
mem[16'h8ED4] = 8'h06;
mem[16'h8ED5] = 8'h00;
mem[16'h8ED6] = 8'h00;
mem[16'h8ED7] = 8'h00;
mem[16'h8ED8] = 8'h00;
mem[16'h8ED9] = 8'h00;
mem[16'h8EDA] = 8'h00;
mem[16'h8EDB] = 8'h00;
mem[16'h8EDC] = 8'h00;
mem[16'h8EDD] = 8'h80;
mem[16'h8EDE] = 8'h80;
mem[16'h8EDF] = 8'h80;
mem[16'h8EE0] = 8'h80;
mem[16'h8EE1] = 8'h80;
mem[16'h8EE2] = 8'h80;
mem[16'h8EE3] = 8'h80;
mem[16'h8EE4] = 8'h80;
mem[16'h8EE5] = 8'h00;
mem[16'h8EE6] = 8'h00;
mem[16'h8EE7] = 8'h00;
mem[16'h8EE8] = 8'h00;
mem[16'h8EE9] = 8'h00;
mem[16'h8EEA] = 8'h00;
mem[16'h8EEB] = 8'h00;
mem[16'h8EEC] = 8'h00;
mem[16'h8EED] = 8'h80;
mem[16'h8EEE] = 8'h80;
mem[16'h8EEF] = 8'h80;
mem[16'h8EF0] = 8'h80;
mem[16'h8EF1] = 8'h80;
mem[16'h8EF2] = 8'h80;
mem[16'h8EF3] = 8'h80;
mem[16'h8EF4] = 8'h80;
mem[16'h8EF5] = 8'h00;
mem[16'h8EF6] = 8'h00;
mem[16'h8EF7] = 8'h00;
mem[16'h8EF8] = 8'h00;
mem[16'h8EF9] = 8'h00;
mem[16'h8EFA] = 8'h00;
mem[16'h8EFB] = 8'h00;
mem[16'h8EFC] = 8'h00;
mem[16'h8EFD] = 8'h80;
mem[16'h8EFE] = 8'h80;
mem[16'h8EFF] = 8'h80;
mem[16'h8F00] = 8'h80;
mem[16'h8F01] = 8'h80;
mem[16'h8F02] = 8'h80;
mem[16'h8F03] = 8'h80;
mem[16'h8F04] = 8'h80;
mem[16'h8F05] = 8'h00;
mem[16'h8F06] = 8'h00;
mem[16'h8F07] = 8'h00;
mem[16'h8F08] = 8'h00;
mem[16'h8F09] = 8'h00;
mem[16'h8F0A] = 8'h00;
mem[16'h8F0B] = 8'h00;
mem[16'h8F0C] = 8'h00;
mem[16'h8F0D] = 8'h80;
mem[16'h8F0E] = 8'h80;
mem[16'h8F0F] = 8'h80;
mem[16'h8F10] = 8'h80;
mem[16'h8F11] = 8'h80;
mem[16'h8F12] = 8'h80;
mem[16'h8F13] = 8'h80;
mem[16'h8F14] = 8'h80;
mem[16'h8F15] = 8'h28;
mem[16'h8F16] = 8'h28;
mem[16'h8F17] = 8'h28;
mem[16'h8F18] = 8'h28;
mem[16'h8F19] = 8'h28;
mem[16'h8F1A] = 8'h28;
mem[16'h8F1B] = 8'h28;
mem[16'h8F1C] = 8'h28;
mem[16'h8F1D] = 8'hA8;
mem[16'h8F1E] = 8'hA8;
mem[16'h8F1F] = 8'hA8;
mem[16'h8F20] = 8'hA8;
mem[16'h8F21] = 8'hA8;
mem[16'h8F22] = 8'hA8;
mem[16'h8F23] = 8'hA8;
mem[16'h8F24] = 8'hA8;
mem[16'h8F25] = 8'h28;
mem[16'h8F26] = 8'h28;
mem[16'h8F27] = 8'h28;
mem[16'h8F28] = 8'h28;
mem[16'h8F29] = 8'h28;
mem[16'h8F2A] = 8'h28;
mem[16'h8F2B] = 8'h28;
mem[16'h8F2C] = 8'h28;
mem[16'h8F2D] = 8'hA8;
mem[16'h8F2E] = 8'hA8;
mem[16'h8F2F] = 8'hA8;
mem[16'h8F30] = 8'hA8;
mem[16'h8F31] = 8'hA8;
mem[16'h8F32] = 8'hA8;
mem[16'h8F33] = 8'hA8;
mem[16'h8F34] = 8'hA8;
mem[16'h8F35] = 8'h28;
mem[16'h8F36] = 8'h28;
mem[16'h8F37] = 8'h28;
mem[16'h8F38] = 8'h28;
mem[16'h8F39] = 8'h28;
mem[16'h8F3A] = 8'h28;
mem[16'h8F3B] = 8'h28;
mem[16'h8F3C] = 8'h28;
mem[16'h8F3D] = 8'hA8;
mem[16'h8F3E] = 8'hA8;
mem[16'h8F3F] = 8'hA8;
mem[16'h8F40] = 8'hA8;
mem[16'h8F41] = 8'hA8;
mem[16'h8F42] = 8'hA8;
mem[16'h8F43] = 8'hA8;
mem[16'h8F44] = 8'hA8;
mem[16'h8F45] = 8'h28;
mem[16'h8F46] = 8'h28;
mem[16'h8F47] = 8'h28;
mem[16'h8F48] = 8'h28;
mem[16'h8F49] = 8'h28;
mem[16'h8F4A] = 8'h28;
mem[16'h8F4B] = 8'h28;
mem[16'h8F4C] = 8'h28;
mem[16'h8F4D] = 8'hA8;
mem[16'h8F4E] = 8'hA8;
mem[16'h8F4F] = 8'hA8;
mem[16'h8F50] = 8'hA8;
mem[16'h8F51] = 8'hA8;
mem[16'h8F52] = 8'hA8;
mem[16'h8F53] = 8'hA8;
mem[16'h8F54] = 8'hA8;
mem[16'h8F55] = 8'h50;
mem[16'h8F56] = 8'h50;
mem[16'h8F57] = 8'h50;
mem[16'h8F58] = 8'h50;
mem[16'h8F59] = 8'h50;
mem[16'h8F5A] = 8'h50;
mem[16'h8F5B] = 8'h50;
mem[16'h8F5C] = 8'h50;
mem[16'h8F5D] = 8'hD0;
mem[16'h8F5E] = 8'hD0;
mem[16'h8F5F] = 8'hD0;
mem[16'h8F60] = 8'hD0;
mem[16'h8F61] = 8'hD0;
mem[16'h8F62] = 8'hD0;
mem[16'h8F63] = 8'hD0;
mem[16'h8F64] = 8'hD0;
mem[16'h8F65] = 8'h50;
mem[16'h8F66] = 8'h50;
mem[16'h8F67] = 8'h50;
mem[16'h8F68] = 8'h50;
mem[16'h8F69] = 8'h50;
mem[16'h8F6A] = 8'h50;
mem[16'h8F6B] = 8'h50;
mem[16'h8F6C] = 8'h50;
mem[16'h8F6D] = 8'hD0;
mem[16'h8F6E] = 8'hD0;
mem[16'h8F6F] = 8'hD0;
mem[16'h8F70] = 8'hD0;
mem[16'h8F71] = 8'hD0;
mem[16'h8F72] = 8'hD0;
mem[16'h8F73] = 8'hD0;
mem[16'h8F74] = 8'hD0;
mem[16'h8F75] = 8'h50;
mem[16'h8F76] = 8'h50;
mem[16'h8F77] = 8'h50;
mem[16'h8F78] = 8'h50;
mem[16'h8F79] = 8'h50;
mem[16'h8F7A] = 8'h50;
mem[16'h8F7B] = 8'h50;
mem[16'h8F7C] = 8'h50;
mem[16'h8F7D] = 8'hD0;
mem[16'h8F7E] = 8'hD0;
mem[16'h8F7F] = 8'hD0;
mem[16'h8F80] = 8'hD0;
mem[16'h8F81] = 8'hD0;
mem[16'h8F82] = 8'hD0;
mem[16'h8F83] = 8'hD0;
mem[16'h8F84] = 8'hD0;
mem[16'h8F85] = 8'h50;
mem[16'h8F86] = 8'h50;
mem[16'h8F87] = 8'h50;
mem[16'h8F88] = 8'h50;
mem[16'h8F89] = 8'h50;
mem[16'h8F8A] = 8'h50;
mem[16'h8F8B] = 8'h50;
mem[16'h8F8C] = 8'h50;
mem[16'h8F8D] = 8'hD0;
mem[16'h8F8E] = 8'hD0;
mem[16'h8F8F] = 8'hD0;
mem[16'h8F90] = 8'hD0;
mem[16'h8F91] = 8'hD0;
mem[16'h8F92] = 8'hD0;
mem[16'h8F93] = 8'hD0;
mem[16'h8F94] = 8'hD0;
mem[16'h8F95] = 8'h20;
mem[16'h8F96] = 8'h24;
mem[16'h8F97] = 8'h28;
mem[16'h8F98] = 8'h2C;
mem[16'h8F99] = 8'h30;
mem[16'h8F9A] = 8'h34;
mem[16'h8F9B] = 8'h38;
mem[16'h8F9C] = 8'h3C;
mem[16'h8F9D] = 8'h20;
mem[16'h8F9E] = 8'h24;
mem[16'h8F9F] = 8'h28;
mem[16'h8FA0] = 8'h2C;
mem[16'h8FA1] = 8'h30;
mem[16'h8FA2] = 8'h34;
mem[16'h8FA3] = 8'h38;
mem[16'h8FA4] = 8'h3C;
mem[16'h8FA5] = 8'h21;
mem[16'h8FA6] = 8'h25;
mem[16'h8FA7] = 8'h29;
mem[16'h8FA8] = 8'h2D;
mem[16'h8FA9] = 8'h31;
mem[16'h8FAA] = 8'h35;
mem[16'h8FAB] = 8'h39;
mem[16'h8FAC] = 8'h3D;
mem[16'h8FAD] = 8'h21;
mem[16'h8FAE] = 8'h25;
mem[16'h8FAF] = 8'h29;
mem[16'h8FB0] = 8'h2D;
mem[16'h8FB1] = 8'h31;
mem[16'h8FB2] = 8'h35;
mem[16'h8FB3] = 8'h39;
mem[16'h8FB4] = 8'h3D;
mem[16'h8FB5] = 8'h22;
mem[16'h8FB6] = 8'h26;
mem[16'h8FB7] = 8'h2A;
mem[16'h8FB8] = 8'h2E;
mem[16'h8FB9] = 8'h32;
mem[16'h8FBA] = 8'h36;
mem[16'h8FBB] = 8'h3A;
mem[16'h8FBC] = 8'h3E;
mem[16'h8FBD] = 8'h22;
mem[16'h8FBE] = 8'h26;
mem[16'h8FBF] = 8'h2A;
mem[16'h8FC0] = 8'h2E;
mem[16'h8FC1] = 8'h32;
mem[16'h8FC2] = 8'h36;
mem[16'h8FC3] = 8'h3A;
mem[16'h8FC4] = 8'h3E;
mem[16'h8FC5] = 8'h23;
mem[16'h8FC6] = 8'h27;
mem[16'h8FC7] = 8'h2B;
mem[16'h8FC8] = 8'h2F;
mem[16'h8FC9] = 8'h33;
mem[16'h8FCA] = 8'h37;
mem[16'h8FCB] = 8'h3B;
mem[16'h8FCC] = 8'h3F;
mem[16'h8FCD] = 8'h23;
mem[16'h8FCE] = 8'h27;
mem[16'h8FCF] = 8'h2B;
mem[16'h8FD0] = 8'h2F;
mem[16'h8FD1] = 8'h33;
mem[16'h8FD2] = 8'h37;
mem[16'h8FD3] = 8'h3B;
mem[16'h8FD4] = 8'h3F;
mem[16'h8FD5] = 8'h20;
mem[16'h8FD6] = 8'h24;
mem[16'h8FD7] = 8'h28;
mem[16'h8FD8] = 8'h2C;
mem[16'h8FD9] = 8'h30;
mem[16'h8FDA] = 8'h34;
mem[16'h8FDB] = 8'h38;
mem[16'h8FDC] = 8'h3C;
mem[16'h8FDD] = 8'h20;
mem[16'h8FDE] = 8'h24;
mem[16'h8FDF] = 8'h28;
mem[16'h8FE0] = 8'h2C;
mem[16'h8FE1] = 8'h30;
mem[16'h8FE2] = 8'h34;
mem[16'h8FE3] = 8'h38;
mem[16'h8FE4] = 8'h3C;
mem[16'h8FE5] = 8'h21;
mem[16'h8FE6] = 8'h25;
mem[16'h8FE7] = 8'h29;
mem[16'h8FE8] = 8'h2D;
mem[16'h8FE9] = 8'h31;
mem[16'h8FEA] = 8'h35;
mem[16'h8FEB] = 8'h39;
mem[16'h8FEC] = 8'h3D;
mem[16'h8FED] = 8'h21;
mem[16'h8FEE] = 8'h25;
mem[16'h8FEF] = 8'h29;
mem[16'h8FF0] = 8'h2D;
mem[16'h8FF1] = 8'h31;
mem[16'h8FF2] = 8'h35;
mem[16'h8FF3] = 8'h39;
mem[16'h8FF4] = 8'h3D;
mem[16'h8FF5] = 8'h22;
mem[16'h8FF6] = 8'h26;
mem[16'h8FF7] = 8'h2A;
mem[16'h8FF8] = 8'h2E;
mem[16'h8FF9] = 8'h32;
mem[16'h8FFA] = 8'h36;
mem[16'h8FFB] = 8'h3A;
mem[16'h8FFC] = 8'h3E;
mem[16'h8FFD] = 8'h22;
mem[16'h8FFE] = 8'h26;
mem[16'h8FFF] = 8'h2A;
mem[16'h9000] = 8'h2E;
mem[16'h9001] = 8'h32;
mem[16'h9002] = 8'h36;
mem[16'h9003] = 8'h3A;
mem[16'h9004] = 8'h3E;
mem[16'h9005] = 8'h23;
mem[16'h9006] = 8'h27;
mem[16'h9007] = 8'h2B;
mem[16'h9008] = 8'h2F;
mem[16'h9009] = 8'h33;
mem[16'h900A] = 8'h37;
mem[16'h900B] = 8'h3B;
mem[16'h900C] = 8'h3F;
mem[16'h900D] = 8'h23;
mem[16'h900E] = 8'h27;
mem[16'h900F] = 8'h2B;
mem[16'h9010] = 8'h2F;
mem[16'h9011] = 8'h33;
mem[16'h9012] = 8'h37;
mem[16'h9013] = 8'h3B;
mem[16'h9014] = 8'h3F;
mem[16'h9015] = 8'h20;
mem[16'h9016] = 8'h24;
mem[16'h9017] = 8'h28;
mem[16'h9018] = 8'h2C;
mem[16'h9019] = 8'h30;
mem[16'h901A] = 8'h34;
mem[16'h901B] = 8'h38;
mem[16'h901C] = 8'h3C;
mem[16'h901D] = 8'h20;
mem[16'h901E] = 8'h24;
mem[16'h901F] = 8'h28;
mem[16'h9020] = 8'h2C;
mem[16'h9021] = 8'h30;
mem[16'h9022] = 8'h34;
mem[16'h9023] = 8'h38;
mem[16'h9024] = 8'h3C;
mem[16'h9025] = 8'h21;
mem[16'h9026] = 8'h25;
mem[16'h9027] = 8'h29;
mem[16'h9028] = 8'h2D;
mem[16'h9029] = 8'h31;
mem[16'h902A] = 8'h35;
mem[16'h902B] = 8'h39;
mem[16'h902C] = 8'h3D;
mem[16'h902D] = 8'h21;
mem[16'h902E] = 8'h25;
mem[16'h902F] = 8'h29;
mem[16'h9030] = 8'h2D;
mem[16'h9031] = 8'h31;
mem[16'h9032] = 8'h35;
mem[16'h9033] = 8'h39;
mem[16'h9034] = 8'h3D;
mem[16'h9035] = 8'h22;
mem[16'h9036] = 8'h26;
mem[16'h9037] = 8'h2A;
mem[16'h9038] = 8'h2E;
mem[16'h9039] = 8'h32;
mem[16'h903A] = 8'h36;
mem[16'h903B] = 8'h3A;
mem[16'h903C] = 8'h3E;
mem[16'h903D] = 8'h22;
mem[16'h903E] = 8'h26;
mem[16'h903F] = 8'h2A;
mem[16'h9040] = 8'h2E;
mem[16'h9041] = 8'h32;
mem[16'h9042] = 8'h36;
mem[16'h9043] = 8'h3A;
mem[16'h9044] = 8'h3E;
mem[16'h9045] = 8'h23;
mem[16'h9046] = 8'h27;
mem[16'h9047] = 8'h2B;
mem[16'h9048] = 8'h2F;
mem[16'h9049] = 8'h33;
mem[16'h904A] = 8'h37;
mem[16'h904B] = 8'h3B;
mem[16'h904C] = 8'h3F;
mem[16'h904D] = 8'h23;
mem[16'h904E] = 8'h27;
mem[16'h904F] = 8'h2B;
mem[16'h9050] = 8'h2F;
mem[16'h9051] = 8'h33;
mem[16'h9052] = 8'h37;
mem[16'h9053] = 8'h3B;
mem[16'h9054] = 8'h3F;
mem[16'h9055] = 8'hA9;
mem[16'h9056] = 8'h08;
mem[16'h9057] = 8'h8D;
mem[16'h9058] = 8'hA2;
mem[16'h9059] = 8'h55;
mem[16'h905A] = 8'hA9;
mem[16'h905B] = 8'h01;
mem[16'h905C] = 8'h8D;
mem[16'h905D] = 8'hA1;
mem[16'h905E] = 8'h55;
mem[16'h905F] = 8'h20;
mem[16'h9060] = 8'h51;
mem[16'h9061] = 8'h55;
mem[16'h9062] = 8'hAD;
mem[16'h9063] = 8'hA1;
mem[16'h9064] = 8'h55;
mem[16'h9065] = 8'h18;
mem[16'h9066] = 8'h69;
mem[16'h9067] = 8'h08;
mem[16'h9068] = 8'h8D;
mem[16'h9069] = 8'hA1;
mem[16'h906A] = 8'h55;
mem[16'h906B] = 8'h90;
mem[16'h906C] = 8'hF2;
mem[16'h906D] = 8'hAD;
mem[16'h906E] = 8'hA2;
mem[16'h906F] = 8'h55;
mem[16'h9070] = 8'h18;
mem[16'h9071] = 8'h69;
mem[16'h9072] = 8'h05;
mem[16'h9073] = 8'hC9;
mem[16'h9074] = 8'h13;
mem[16'h9075] = 8'hB0;
mem[16'h9076] = 8'h06;
mem[16'h9077] = 8'h8D;
mem[16'h9078] = 8'hA2;
mem[16'h9079] = 8'h55;
mem[16'h907A] = 8'h4C;
mem[16'h907B] = 8'h5A;
mem[16'h907C] = 8'h90;
mem[16'h907D] = 8'hA9;
mem[16'h907E] = 8'h15;
mem[16'h907F] = 8'h20;
mem[16'h9080] = 8'hB2;
mem[16'h9081] = 8'h54;
mem[16'h9082] = 8'hA9;
mem[16'h9083] = 8'h46;
mem[16'h9084] = 8'h20;
mem[16'h9085] = 8'hB2;
mem[16'h9086] = 8'h54;
mem[16'h9087] = 8'hA9;
mem[16'h9088] = 8'h70;
mem[16'h9089] = 8'h20;
mem[16'h908A] = 8'hB2;
mem[16'h908B] = 8'h54;
mem[16'h908C] = 8'hA9;
mem[16'h908D] = 8'hA1;
mem[16'h908E] = 8'h20;
mem[16'h908F] = 8'hB2;
mem[16'h9090] = 8'h54;
mem[16'h9091] = 8'hA9;
mem[16'h9092] = 8'hCB;
mem[16'h9093] = 8'h20;
mem[16'h9094] = 8'hB2;
mem[16'h9095] = 8'h54;
mem[16'h9096] = 8'h60;
mem[16'h9097] = 8'hAD;
mem[16'h9098] = 8'hE6;
mem[16'h9099] = 8'h48;
mem[16'h909A] = 8'hC9;
mem[16'h909B] = 8'h01;
mem[16'h909C] = 8'hF0;
mem[16'h909D] = 8'h34;
mem[16'h909E] = 8'hA9;
mem[16'h909F] = 8'h02;
mem[16'h90A0] = 8'h85;
mem[16'h90A1] = 8'h56;
mem[16'h90A2] = 8'h20;
mem[16'h90A3] = 8'h54;
mem[16'h90A4] = 8'h8B;
mem[16'h90A5] = 8'hAD;
mem[16'h90A6] = 8'hE6;
mem[16'h90A7] = 8'h48;
mem[16'h90A8] = 8'hC9;
mem[16'h90A9] = 8'h02;
mem[16'h90AA] = 8'hF0;
mem[16'h90AB] = 8'h26;
mem[16'h90AC] = 8'hA9;
mem[16'h90AD] = 8'h10;
mem[16'h90AE] = 8'h85;
mem[16'h90AF] = 8'h56;
mem[16'h90B0] = 8'h20;
mem[16'h90B1] = 8'h54;
mem[16'h90B2] = 8'h8B;
mem[16'h90B3] = 8'hAD;
mem[16'h90B4] = 8'hE6;
mem[16'h90B5] = 8'h48;
mem[16'h90B6] = 8'hC9;
mem[16'h90B7] = 8'h03;
mem[16'h90B8] = 8'hF0;
mem[16'h90B9] = 8'h18;
mem[16'h90BA] = 8'hA9;
mem[16'h90BB] = 8'h1E;
mem[16'h90BC] = 8'h85;
mem[16'h90BD] = 8'h56;
mem[16'h90BE] = 8'h20;
mem[16'h90BF] = 8'h54;
mem[16'h90C0] = 8'h8B;
mem[16'h90C1] = 8'hAD;
mem[16'h90C2] = 8'hE6;
mem[16'h90C3] = 8'h48;
mem[16'h90C4] = 8'hC9;
mem[16'h90C5] = 8'h04;
mem[16'h90C6] = 8'hF0;
mem[16'h90C7] = 8'h0A;
mem[16'h90C8] = 8'hA9;
mem[16'h90C9] = 8'h2C;
mem[16'h90CA] = 8'h85;
mem[16'h90CB] = 8'h56;
mem[16'h90CC] = 8'h8D;
mem[16'h90CD] = 8'hD3;
mem[16'h90CE] = 8'h90;
mem[16'h90CF] = 8'h20;
mem[16'h90D0] = 8'h54;
mem[16'h90D1] = 8'h8B;
mem[16'h90D2] = 8'h60;
mem[16'h90D3] = 8'h2C;
mem[16'h90D4] = 8'hC6;
mem[16'h90D5] = 8'h73;
mem[16'h90D6] = 8'hF0;
mem[16'h90D7] = 8'h03;
mem[16'h90D8] = 8'h4C;
mem[16'h90D9] = 8'h10;
mem[16'h90DA] = 8'h91;
mem[16'h90DB] = 8'hAD;
mem[16'h90DC] = 8'hE0;
mem[16'h90DD] = 8'h91;
mem[16'h90DE] = 8'h85;
mem[16'h90DF] = 8'h73;
mem[16'h90E0] = 8'hF8;
mem[16'h90E1] = 8'hA5;
mem[16'h90E2] = 8'h74;
mem[16'h90E3] = 8'h38;
mem[16'h90E4] = 8'hE9;
mem[16'h90E5] = 8'h01;
mem[16'h90E6] = 8'h85;
mem[16'h90E7] = 8'h74;
mem[16'h90E8] = 8'hD8;
mem[16'h90E9] = 8'hEE;
mem[16'h90EA] = 8'hD8;
mem[16'h90EB] = 8'h91;
mem[16'h90EC] = 8'h20;
mem[16'h90ED] = 8'h2D;
mem[16'h90EE] = 8'h92;
mem[16'h90EF] = 8'hA5;
mem[16'h90F0] = 8'h74;
mem[16'h90F1] = 8'hC9;
mem[16'h90F2] = 8'h10;
mem[16'h90F3] = 8'hD0;
mem[16'h90F4] = 8'h05;
mem[16'h90F5] = 8'h20;
mem[16'h90F6] = 8'h56;
mem[16'h90F7] = 8'h92;
mem[16'h90F8] = 8'hA5;
mem[16'h90F9] = 8'h74;
mem[16'h90FA] = 8'hC9;
mem[16'h90FB] = 8'h00;
mem[16'h90FC] = 8'hD0;
mem[16'h90FD] = 8'h12;
mem[16'h90FE] = 8'h20;
mem[16'h90FF] = 8'hAE;
mem[16'h9100] = 8'h4C;
mem[16'h9101] = 8'h20;
mem[16'h9102] = 8'hBE;
mem[16'h9103] = 8'h7E;
mem[16'h9104] = 8'h20;
mem[16'h9105] = 8'h6D;
mem[16'h9106] = 8'h4C;
mem[16'h9107] = 8'h20;
mem[16'h9108] = 8'hBE;
mem[16'h9109] = 8'h7E;
mem[16'h910A] = 8'h20;
mem[16'h910B] = 8'hA6;
mem[16'h910C] = 8'h6D;
mem[16'h910D] = 8'h4C;
mem[16'h910E] = 8'h97;
mem[16'h910F] = 8'h48;
mem[16'h9110] = 8'hCE;
mem[16'h9111] = 8'hDC;
mem[16'h9112] = 8'h91;
mem[16'h9113] = 8'hD0;
mem[16'h9114] = 8'h7E;
mem[16'h9115] = 8'hA9;
mem[16'h9116] = 8'h01;
mem[16'h9117] = 8'h8D;
mem[16'h9118] = 8'hDC;
mem[16'h9119] = 8'h91;
mem[16'h911A] = 8'hAD;
mem[16'h911B] = 8'h13;
mem[16'h911C] = 8'h87;
mem[16'h911D] = 8'h29;
mem[16'h911E] = 8'h0F;
mem[16'h911F] = 8'h8D;
mem[16'h9120] = 8'hC5;
mem[16'h9121] = 8'h5E;
mem[16'h9122] = 8'hCD;
mem[16'h9123] = 8'hAF;
mem[16'h9124] = 8'h4A;
mem[16'h9125] = 8'hB0;
mem[16'h9126] = 8'h1D;
mem[16'h9127] = 8'hA9;
mem[16'h9128] = 8'h00;
mem[16'h9129] = 8'h18;
mem[16'h912A] = 8'h6D;
mem[16'h912B] = 8'h63;
mem[16'h912C] = 8'h5E;
mem[16'h912D] = 8'hCD;
mem[16'h912E] = 8'hC5;
mem[16'h912F] = 8'h5E;
mem[16'h9130] = 8'hB0;
mem[16'h9131] = 8'h08;
mem[16'h9132] = 8'hCD;
mem[16'h9133] = 8'hAF;
mem[16'h9134] = 8'h4A;
mem[16'h9135] = 8'h90;
mem[16'h9136] = 8'hF2;
mem[16'h9137] = 8'h4C;
mem[16'h9138] = 8'h44;
mem[16'h9139] = 8'h91;
mem[16'h913A] = 8'h8D;
mem[16'h913B] = 8'hC5;
mem[16'h913C] = 8'h5E;
mem[16'h913D] = 8'h38;
mem[16'h913E] = 8'hED;
mem[16'h913F] = 8'h63;
mem[16'h9140] = 8'h5E;
mem[16'h9141] = 8'h4C;
mem[16'h9142] = 8'h66;
mem[16'h9143] = 8'h91;
mem[16'h9144] = 8'hAD;
mem[16'h9145] = 8'hC5;
mem[16'h9146] = 8'h5E;
mem[16'h9147] = 8'hCD;
mem[16'h9148] = 8'hB0;
mem[16'h9149] = 8'h4A;
mem[16'h914A] = 8'hB0;
mem[16'h914B] = 8'h47;
mem[16'h914C] = 8'hA9;
mem[16'h914D] = 8'h08;
mem[16'h914E] = 8'h18;
mem[16'h914F] = 8'h6D;
mem[16'h9150] = 8'hC4;
mem[16'h9151] = 8'h5E;
mem[16'h9152] = 8'hCD;
mem[16'h9153] = 8'hC5;
mem[16'h9154] = 8'h5E;
mem[16'h9155] = 8'hB0;
mem[16'h9156] = 8'h08;
mem[16'h9157] = 8'hCD;
mem[16'h9158] = 8'hB0;
mem[16'h9159] = 8'h4A;
mem[16'h915A] = 8'h90;
mem[16'h915B] = 8'hF2;
mem[16'h915C] = 8'h4C;
mem[16'h915D] = 8'h93;
mem[16'h915E] = 8'h91;
mem[16'h915F] = 8'h8D;
mem[16'h9160] = 8'hC5;
mem[16'h9161] = 8'h5E;
mem[16'h9162] = 8'h38;
mem[16'h9163] = 8'hED;
mem[16'h9164] = 8'hC4;
mem[16'h9165] = 8'h5E;
mem[16'h9166] = 8'hAA;
mem[16'h9167] = 8'hBD;
mem[16'h9168] = 8'h83;
mem[16'h9169] = 8'h5B;
mem[16'h916A] = 8'hC9;
mem[16'h916B] = 8'h0D;
mem[16'h916C] = 8'h90;
mem[16'h916D] = 8'h25;
mem[16'h916E] = 8'hC9;
mem[16'h916F] = 8'h14;
mem[16'h9170] = 8'hB0;
mem[16'h9171] = 8'h21;
mem[16'h9172] = 8'hBD;
mem[16'h9173] = 8'h75;
mem[16'h9174] = 8'h5B;
mem[16'h9175] = 8'hD0;
mem[16'h9176] = 8'h1C;
mem[16'h9177] = 8'hBD;
mem[16'h9178] = 8'h2C;
mem[16'h9179] = 8'h5F;
mem[16'h917A] = 8'hC9;
mem[16'h917B] = 8'h0A;
mem[16'h917C] = 8'h90;
mem[16'h917D] = 8'h15;
mem[16'h917E] = 8'hC9;
mem[16'h917F] = 8'hFA;
mem[16'h9180] = 8'hB0;
mem[16'h9181] = 8'h11;
mem[16'h9182] = 8'hAD;
mem[16'h9183] = 8'hDD;
mem[16'h9184] = 8'h91;
mem[16'h9185] = 8'h8D;
mem[16'h9186] = 8'hDC;
mem[16'h9187] = 8'h91;
mem[16'h9188] = 8'hA9;
mem[16'h9189] = 8'h24;
mem[16'h918A] = 8'h9D;
mem[16'h918B] = 8'h75;
mem[16'h918C] = 8'h5B;
mem[16'h918D] = 8'hE8;
mem[16'h918E] = 8'hEC;
mem[16'h918F] = 8'hC5;
mem[16'h9190] = 8'h5E;
mem[16'h9191] = 8'hD0;
mem[16'h9192] = 8'hF7;
mem[16'h9193] = 8'hAD;
mem[16'h9194] = 8'hDA;
mem[16'h9195] = 8'h91;
mem[16'h9196] = 8'hF0;
mem[16'h9197] = 8'h19;
mem[16'h9198] = 8'hCE;
mem[16'h9199] = 8'hDA;
mem[16'h919A] = 8'h91;
mem[16'h919B] = 8'hD0;
mem[16'h919C] = 8'h14;
mem[16'h919D] = 8'hAD;
mem[16'h919E] = 8'hDE;
mem[16'h919F] = 8'h91;
mem[16'h91A0] = 8'h8D;
mem[16'h91A1] = 8'hDA;
mem[16'h91A2] = 8'h91;
mem[16'h91A3] = 8'h20;
mem[16'h91A4] = 8'h61;
mem[16'h91A5] = 8'h77;
mem[16'h91A6] = 8'hAD;
mem[16'h91A7] = 8'hB0;
mem[16'h91A8] = 8'h85;
mem[16'h91A9] = 8'hD0;
mem[16'h91AA] = 8'h06;
mem[16'h91AB] = 8'hAD;
mem[16'h91AC] = 8'hB1;
mem[16'h91AD] = 8'h85;
mem[16'h91AE] = 8'h8D;
mem[16'h91AF] = 8'hB0;
mem[16'h91B0] = 8'h85;
mem[16'h91B1] = 8'hAD;
mem[16'h91B2] = 8'hDB;
mem[16'h91B3] = 8'h91;
mem[16'h91B4] = 8'hF0;
mem[16'h91B5] = 8'h0E;
mem[16'h91B6] = 8'hCE;
mem[16'h91B7] = 8'hDB;
mem[16'h91B8] = 8'h91;
mem[16'h91B9] = 8'hD0;
mem[16'h91BA] = 8'h09;
mem[16'h91BB] = 8'hAD;
mem[16'h91BC] = 8'hDF;
mem[16'h91BD] = 8'h91;
mem[16'h91BE] = 8'h8D;
mem[16'h91BF] = 8'hDB;
mem[16'h91C0] = 8'h91;
mem[16'h91C1] = 8'h20;
mem[16'h91C2] = 8'hB4;
mem[16'h91C3] = 8'h79;
mem[16'h91C4] = 8'hAD;
mem[16'h91C5] = 8'hB0;
mem[16'h91C6] = 8'h85;
mem[16'h91C7] = 8'hF0;
mem[16'h91C8] = 8'h03;
mem[16'h91C9] = 8'hCE;
mem[16'h91CA] = 8'hB0;
mem[16'h91CB] = 8'h85;
mem[16'h91CC] = 8'hAD;
mem[16'h91CD] = 8'hD8;
mem[16'h91CE] = 8'h91;
mem[16'h91CF] = 8'hCD;
mem[16'h91D0] = 8'hD9;
mem[16'h91D1] = 8'h91;
mem[16'h91D2] = 8'hD0;
mem[16'h91D3] = 8'h03;
mem[16'h91D4] = 8'h20;
mem[16'h91D5] = 8'hE1;
mem[16'h91D6] = 8'h91;
mem[16'h91D7] = 8'h60;
mem[16'h91D8] = 8'h1A;
mem[16'h91D9] = 8'hC8;
mem[16'h91DA] = 8'h00;
mem[16'h91DB] = 8'h00;
mem[16'h91DC] = 8'h28;
mem[16'h91DD] = 8'h28;
mem[16'h91DE] = 8'h00;
mem[16'h91DF] = 8'h00;
mem[16'h91E0] = 8'h06;
mem[16'h91E1] = 8'hAD;
mem[16'h91E2] = 8'h13;
mem[16'h91E3] = 8'h87;
mem[16'h91E4] = 8'h8D;
mem[16'h91E5] = 8'hD9;
mem[16'h91E6] = 8'h91;
mem[16'h91E7] = 8'hAD;
mem[16'h91E8] = 8'hB9;
mem[16'h91E9] = 8'h4A;
mem[16'h91EA] = 8'hC9;
mem[16'h91EB] = 8'h03;
mem[16'h91EC] = 8'hF0;
mem[16'h91ED] = 8'h1F;
mem[16'h91EE] = 8'hA9;
mem[16'h91EF] = 8'h01;
mem[16'h91F0] = 8'h8D;
mem[16'h91F1] = 8'hB7;
mem[16'h91F2] = 8'h4A;
mem[16'h91F3] = 8'h8D;
mem[16'h91F4] = 8'hB6;
mem[16'h91F5] = 8'h4A;
mem[16'h91F6] = 8'hA9;
mem[16'h91F7] = 8'h02;
mem[16'h91F8] = 8'h8D;
mem[16'h91F9] = 8'hB4;
mem[16'h91FA] = 8'h4A;
mem[16'h91FB] = 8'h8D;
mem[16'h91FC] = 8'hB5;
mem[16'h91FD] = 8'h4A;
mem[16'h91FE] = 8'h8D;
mem[16'h91FF] = 8'hBA;
mem[16'h9200] = 8'h4A;
mem[16'h9201] = 8'h8D;
mem[16'h9202] = 8'hBB;
mem[16'h9203] = 8'h4A;
mem[16'h9204] = 8'h8D;
mem[16'h9205] = 8'hBC;
mem[16'h9206] = 8'h4A;
mem[16'h9207] = 8'hA9;
mem[16'h9208] = 8'h03;
mem[16'h9209] = 8'h8D;
mem[16'h920A] = 8'hB9;
mem[16'h920B] = 8'h4A;
mem[16'h920C] = 8'h60;
mem[16'h920D] = 8'hA9;
mem[16'h920E] = 8'h01;
mem[16'h920F] = 8'h8D;
mem[16'h9210] = 8'hB4;
mem[16'h9211] = 8'h4A;
mem[16'h9212] = 8'h8D;
mem[16'h9213] = 8'hB5;
mem[16'h9214] = 8'h4A;
mem[16'h9215] = 8'h8D;
mem[16'h9216] = 8'hBA;
mem[16'h9217] = 8'h4A;
mem[16'h9218] = 8'h8D;
mem[16'h9219] = 8'hBB;
mem[16'h921A] = 8'h4A;
mem[16'h921B] = 8'h8D;
mem[16'h921C] = 8'hBC;
mem[16'h921D] = 8'h4A;
mem[16'h921E] = 8'hA9;
mem[16'h921F] = 8'h02;
mem[16'h9220] = 8'h8D;
mem[16'h9221] = 8'hB6;
mem[16'h9222] = 8'h4A;
mem[16'h9223] = 8'h8D;
mem[16'h9224] = 8'hB8;
mem[16'h9225] = 8'h4A;
mem[16'h9226] = 8'h8D;
mem[16'h9227] = 8'hB9;
mem[16'h9228] = 8'h4A;
mem[16'h9229] = 8'h8D;
mem[16'h922A] = 8'hB7;
mem[16'h922B] = 8'h4A;
mem[16'h922C] = 8'h60;
mem[16'h922D] = 8'hAE;
mem[16'h922E] = 8'h34;
mem[16'h922F] = 8'h45;
mem[16'h9230] = 8'hBD;
mem[16'h9231] = 8'hD5;
mem[16'h9232] = 8'h8E;
mem[16'h9233] = 8'h85;
mem[16'h9234] = 8'h59;
mem[16'h9235] = 8'hBD;
mem[16'h9236] = 8'h95;
mem[16'h9237] = 8'h8F;
mem[16'h9238] = 8'h85;
mem[16'h9239] = 8'h5A;
mem[16'h923A] = 8'hA0;
mem[16'h923B] = 8'h27;
mem[16'h923C] = 8'hA9;
mem[16'h923D] = 8'h00;
mem[16'h923E] = 8'h91;
mem[16'h923F] = 8'h59;
mem[16'h9240] = 8'hEE;
mem[16'h9241] = 8'h34;
mem[16'h9242] = 8'h45;
mem[16'h9243] = 8'hE8;
mem[16'h9244] = 8'hBD;
mem[16'h9245] = 8'hD5;
mem[16'h9246] = 8'h8E;
mem[16'h9247] = 8'h85;
mem[16'h9248] = 8'h59;
mem[16'h9249] = 8'hBD;
mem[16'h924A] = 8'h95;
mem[16'h924B] = 8'h8F;
mem[16'h924C] = 8'h85;
mem[16'h924D] = 8'h5A;
mem[16'h924E] = 8'hA9;
mem[16'h924F] = 8'h00;
mem[16'h9250] = 8'h91;
mem[16'h9251] = 8'h59;
mem[16'h9252] = 8'hEE;
mem[16'h9253] = 8'h34;
mem[16'h9254] = 8'h45;
mem[16'h9255] = 8'h60;
mem[16'h9256] = 8'hAE;
mem[16'h9257] = 8'h34;
mem[16'h9258] = 8'h45;
mem[16'h9259] = 8'hBD;
mem[16'h925A] = 8'hD5;
mem[16'h925B] = 8'h8E;
mem[16'h925C] = 8'h85;
mem[16'h925D] = 8'h59;
mem[16'h925E] = 8'hBD;
mem[16'h925F] = 8'h95;
mem[16'h9260] = 8'h8F;
mem[16'h9261] = 8'h85;
mem[16'h9262] = 8'h5A;
mem[16'h9263] = 8'hA0;
mem[16'h9264] = 8'h27;
mem[16'h9265] = 8'hB1;
mem[16'h9266] = 8'h59;
mem[16'h9267] = 8'h09;
mem[16'h9268] = 8'h80;
mem[16'h9269] = 8'h91;
mem[16'h926A] = 8'h59;
mem[16'h926B] = 8'hE8;
mem[16'h926C] = 8'hE0;
mem[16'h926D] = 8'hBE;
mem[16'h926E] = 8'hD0;
mem[16'h926F] = 8'hE9;
mem[16'h9270] = 8'h20;
mem[16'h9271] = 8'h74;
mem[16'h9272] = 8'h92;
mem[16'h9273] = 8'h60;
mem[16'h9274] = 8'hA9;
mem[16'h9275] = 8'h00;
mem[16'h9276] = 8'h85;
mem[16'h9277] = 8'h55;
mem[16'h9278] = 8'hA9;
mem[16'h9279] = 8'h06;
mem[16'h927A] = 8'h85;
mem[16'h927B] = 8'h52;
mem[16'h927C] = 8'h85;
mem[16'h927D] = 8'h53;
mem[16'h927E] = 8'hAD;
mem[16'h927F] = 8'hB1;
mem[16'h9280] = 8'h92;
mem[16'h9281] = 8'h85;
mem[16'h9282] = 8'h50;
mem[16'h9283] = 8'h20;
mem[16'h9284] = 8'h00;
mem[16'h9285] = 8'h65;
mem[16'h9286] = 8'hA9;
mem[16'h9287] = 8'h06;
mem[16'h9288] = 8'h85;
mem[16'h9289] = 8'h52;
mem[16'h928A] = 8'h85;
mem[16'h928B] = 8'h53;
mem[16'h928C] = 8'hAD;
mem[16'h928D] = 8'hB2;
mem[16'h928E] = 8'h92;
mem[16'h928F] = 8'h85;
mem[16'h9290] = 8'h50;
mem[16'h9291] = 8'h20;
mem[16'h9292] = 8'h00;
mem[16'h9293] = 8'h65;
mem[16'h9294] = 8'hA9;
mem[16'h9295] = 8'h06;
mem[16'h9296] = 8'h85;
mem[16'h9297] = 8'h52;
mem[16'h9298] = 8'h85;
mem[16'h9299] = 8'h53;
mem[16'h929A] = 8'hAD;
mem[16'h929B] = 8'hB3;
mem[16'h929C] = 8'h92;
mem[16'h929D] = 8'h85;
mem[16'h929E] = 8'h50;
mem[16'h929F] = 8'h20;
mem[16'h92A0] = 8'h00;
mem[16'h92A1] = 8'h65;
mem[16'h92A2] = 8'hA9;
mem[16'h92A3] = 8'h06;
mem[16'h92A4] = 8'h85;
mem[16'h92A5] = 8'h52;
mem[16'h92A6] = 8'h85;
mem[16'h92A7] = 8'h53;
mem[16'h92A8] = 8'hAD;
mem[16'h92A9] = 8'hB4;
mem[16'h92AA] = 8'h92;
mem[16'h92AB] = 8'h85;
mem[16'h92AC] = 8'h50;
mem[16'h92AD] = 8'h20;
mem[16'h92AE] = 8'h00;
mem[16'h92AF] = 8'h65;
mem[16'h92B0] = 8'h60;
mem[16'h92B1] = 8'h22;
mem[16'h92B2] = 8'h2D;
mem[16'h92B3] = 8'h1B;
mem[16'h92B4] = 8'h28;
mem[16'h92B5] = 8'h00;
mem[16'h92B6] = 8'h10;
mem[16'h92B7] = 8'h00;
mem[16'h92B8] = 8'h00;
mem[16'h92B9] = 8'h00;
mem[16'h92BA] = 8'h50;
mem[16'h92BB] = 8'h08;
mem[16'h92BC] = 8'h00;
mem[16'h92BD] = 8'h00;
mem[16'h92BE] = 8'h30;
mem[16'h92BF] = 8'h24;
mem[16'h92C0] = 8'h00;
mem[16'h92C1] = 8'h00;
mem[16'h92C2] = 8'h06;
mem[16'h92C3] = 8'h30;
mem[16'h92C4] = 8'h00;
mem[16'h92C5] = 8'h40;
mem[16'h92C6] = 8'h38;
mem[16'h92C7] = 8'h40;
mem[16'h92C8] = 8'h01;
mem[16'h92C9] = 8'h40;
mem[16'h92CA] = 8'h38;
mem[16'h92CB] = 8'h40;
mem[16'h92CC] = 8'h01;
mem[16'h92CD] = 8'h40;
mem[16'h92CE] = 8'h38;
mem[16'h92CF] = 8'h40;
mem[16'h92D0] = 8'h01;
mem[16'h92D1] = 8'h00;
mem[16'h92D2] = 8'h06;
mem[16'h92D3] = 8'h30;
mem[16'h92D4] = 8'h00;
mem[16'h92D5] = 8'h00;
mem[16'h92D6] = 8'h30;
mem[16'h92D7] = 8'h24;
mem[16'h92D8] = 8'h00;
mem[16'h92D9] = 8'h00;
mem[16'h92DA] = 8'h50;
mem[16'h92DB] = 8'h08;
mem[16'h92DC] = 8'h00;
mem[16'h92DD] = 8'h00;
mem[16'h92DE] = 8'h10;
mem[16'h92DF] = 8'h00;
mem[16'h92E0] = 8'h00;
mem[16'h92E1] = 8'h00;
mem[16'h92E2] = 8'h08;
mem[16'h92E3] = 8'h00;
mem[16'h92E4] = 8'h00;
mem[16'h92E5] = 8'h00;
mem[16'h92E6] = 8'h28;
mem[16'h92E7] = 8'h04;
mem[16'h92E8] = 8'h00;
mem[16'h92E9] = 8'h00;
mem[16'h92EA] = 8'h18;
mem[16'h92EB] = 8'h12;
mem[16'h92EC] = 8'h00;
mem[16'h92ED] = 8'h00;
mem[16'h92EE] = 8'h03;
mem[16'h92EF] = 8'h18;
mem[16'h92F0] = 8'h00;
mem[16'h92F1] = 8'h20;
mem[16'h92F2] = 8'h1C;
mem[16'h92F3] = 8'h60;
mem[16'h92F4] = 8'h00;
mem[16'h92F5] = 8'h20;
mem[16'h92F6] = 8'h1C;
mem[16'h92F7] = 8'h60;
mem[16'h92F8] = 8'h00;
mem[16'h92F9] = 8'h20;
mem[16'h92FA] = 8'h1C;
mem[16'h92FB] = 8'h60;
mem[16'h92FC] = 8'h00;
mem[16'h92FD] = 8'h00;
mem[16'h92FE] = 8'h03;
mem[16'h92FF] = 8'h18;
mem[16'h9300] = 8'h00;
mem[16'h9301] = 8'h00;
mem[16'h9302] = 8'h18;
mem[16'h9303] = 8'h12;
mem[16'h9304] = 8'h00;
mem[16'h9305] = 8'h00;
mem[16'h9306] = 8'h28;
mem[16'h9307] = 8'h04;
mem[16'h9308] = 8'h00;
mem[16'h9309] = 8'h00;
mem[16'h930A] = 8'h08;
mem[16'h930B] = 8'h00;
mem[16'h930C] = 8'h00;
mem[16'h930D] = 8'h00;
mem[16'h930E] = 8'h04;
mem[16'h930F] = 8'h00;
mem[16'h9310] = 8'h00;
mem[16'h9311] = 8'h00;
mem[16'h9312] = 8'h14;
mem[16'h9313] = 8'h02;
mem[16'h9314] = 8'h00;
mem[16'h9315] = 8'h00;
mem[16'h9316] = 8'h0C;
mem[16'h9317] = 8'h09;
mem[16'h9318] = 8'h00;
mem[16'h9319] = 8'h40;
mem[16'h931A] = 8'h01;
mem[16'h931B] = 8'h0C;
mem[16'h931C] = 8'h00;
mem[16'h931D] = 8'h10;
mem[16'h931E] = 8'h0E;
mem[16'h931F] = 8'h30;
mem[16'h9320] = 8'h00;
mem[16'h9321] = 8'h10;
mem[16'h9322] = 8'h0E;
mem[16'h9323] = 8'h30;
mem[16'h9324] = 8'h00;
mem[16'h9325] = 8'h10;
mem[16'h9326] = 8'h0E;
mem[16'h9327] = 8'h30;
mem[16'h9328] = 8'h00;
mem[16'h9329] = 8'h40;
mem[16'h932A] = 8'h01;
mem[16'h932B] = 8'h0C;
mem[16'h932C] = 8'h00;
mem[16'h932D] = 8'h00;
mem[16'h932E] = 8'h0C;
mem[16'h932F] = 8'h09;
mem[16'h9330] = 8'h00;
mem[16'h9331] = 8'h00;
mem[16'h9332] = 8'h14;
mem[16'h9333] = 8'h02;
mem[16'h9334] = 8'h00;
mem[16'h9335] = 8'h00;
mem[16'h9336] = 8'h04;
mem[16'h9337] = 8'h00;
mem[16'h9338] = 8'h00;
mem[16'h9339] = 8'h00;
mem[16'h933A] = 8'h02;
mem[16'h933B] = 8'h00;
mem[16'h933C] = 8'h00;
mem[16'h933D] = 8'h00;
mem[16'h933E] = 8'h0A;
mem[16'h933F] = 8'h01;
mem[16'h9340] = 8'h00;
mem[16'h9341] = 8'h00;
mem[16'h9342] = 8'h46;
mem[16'h9343] = 8'h04;
mem[16'h9344] = 8'h00;
mem[16'h9345] = 8'h60;
mem[16'h9346] = 8'h00;
mem[16'h9347] = 8'h06;
mem[16'h9348] = 8'h00;
mem[16'h9349] = 8'h08;
mem[16'h934A] = 8'h07;
mem[16'h934B] = 8'h18;
mem[16'h934C] = 8'h00;
mem[16'h934D] = 8'h08;
mem[16'h934E] = 8'h07;
mem[16'h934F] = 8'h18;
mem[16'h9350] = 8'h00;
mem[16'h9351] = 8'h08;
mem[16'h9352] = 8'h07;
mem[16'h9353] = 8'h18;
mem[16'h9354] = 8'h00;
mem[16'h9355] = 8'h60;
mem[16'h9356] = 8'h00;
mem[16'h9357] = 8'h06;
mem[16'h9358] = 8'h00;
mem[16'h9359] = 8'h00;
mem[16'h935A] = 8'h46;
mem[16'h935B] = 8'h04;
mem[16'h935C] = 8'h00;
mem[16'h935D] = 8'h00;
mem[16'h935E] = 8'h0A;
mem[16'h935F] = 8'h01;
mem[16'h9360] = 8'h00;
mem[16'h9361] = 8'h00;
mem[16'h9362] = 8'h02;
mem[16'h9363] = 8'h00;
mem[16'h9364] = 8'h00;
mem[16'h9365] = 8'h00;
mem[16'h9366] = 8'h01;
mem[16'h9367] = 8'h00;
mem[16'h9368] = 8'h00;
mem[16'h9369] = 8'h00;
mem[16'h936A] = 8'h45;
mem[16'h936B] = 8'h00;
mem[16'h936C] = 8'h00;
mem[16'h936D] = 8'h00;
mem[16'h936E] = 8'h23;
mem[16'h936F] = 8'h02;
mem[16'h9370] = 8'h00;
mem[16'h9371] = 8'h30;
mem[16'h9372] = 8'h00;
mem[16'h9373] = 8'h03;
mem[16'h9374] = 8'h00;
mem[16'h9375] = 8'h44;
mem[16'h9376] = 8'h03;
mem[16'h9377] = 8'h0C;
mem[16'h9378] = 8'h00;
mem[16'h9379] = 8'h44;
mem[16'h937A] = 8'h03;
mem[16'h937B] = 8'h0C;
mem[16'h937C] = 8'h00;
mem[16'h937D] = 8'h44;
mem[16'h937E] = 8'h03;
mem[16'h937F] = 8'h0C;
mem[16'h9380] = 8'h00;
mem[16'h9381] = 8'h30;
mem[16'h9382] = 8'h00;
mem[16'h9383] = 8'h03;
mem[16'h9384] = 8'h00;
mem[16'h9385] = 8'h00;
mem[16'h9386] = 8'h23;
mem[16'h9387] = 8'h02;
mem[16'h9388] = 8'h00;
mem[16'h9389] = 8'h00;
mem[16'h938A] = 8'h45;
mem[16'h938B] = 8'h00;
mem[16'h938C] = 8'h00;
mem[16'h938D] = 8'h00;
mem[16'h938E] = 8'h01;
mem[16'h938F] = 8'h00;
mem[16'h9390] = 8'h00;
mem[16'h9391] = 8'h40;
mem[16'h9392] = 8'h00;
mem[16'h9393] = 8'h00;
mem[16'h9394] = 8'h00;
mem[16'h9395] = 8'h40;
mem[16'h9396] = 8'h22;
mem[16'h9397] = 8'h00;
mem[16'h9398] = 8'h00;
mem[16'h9399] = 8'h40;
mem[16'h939A] = 8'h11;
mem[16'h939B] = 8'h01;
mem[16'h939C] = 8'h00;
mem[16'h939D] = 8'h18;
mem[16'h939E] = 8'h40;
mem[16'h939F] = 8'h01;
mem[16'h93A0] = 8'h00;
mem[16'h93A1] = 8'h62;
mem[16'h93A2] = 8'h01;
mem[16'h93A3] = 8'h06;
mem[16'h93A4] = 8'h00;
mem[16'h93A5] = 8'h62;
mem[16'h93A6] = 8'h01;
mem[16'h93A7] = 8'h06;
mem[16'h93A8] = 8'h00;
mem[16'h93A9] = 8'h62;
mem[16'h93AA] = 8'h01;
mem[16'h93AB] = 8'h06;
mem[16'h93AC] = 8'h00;
mem[16'h93AD] = 8'h18;
mem[16'h93AE] = 8'h40;
mem[16'h93AF] = 8'h01;
mem[16'h93B0] = 8'h00;
mem[16'h93B1] = 8'h40;
mem[16'h93B2] = 8'h11;
mem[16'h93B3] = 8'h01;
mem[16'h93B4] = 8'h00;
mem[16'h93B5] = 8'h40;
mem[16'h93B6] = 8'h22;
mem[16'h93B7] = 8'h00;
mem[16'h93B8] = 8'h00;
mem[16'h93B9] = 8'h40;
mem[16'h93BA] = 8'h00;
mem[16'h93BB] = 8'h00;
mem[16'h93BC] = 8'h00;
mem[16'h93BD] = 8'h20;
mem[16'h93BE] = 8'h00;
mem[16'h93BF] = 8'h00;
mem[16'h93C0] = 8'h00;
mem[16'h93C1] = 8'h20;
mem[16'h93C2] = 8'h11;
mem[16'h93C3] = 8'h00;
mem[16'h93C4] = 8'h00;
mem[16'h93C5] = 8'h60;
mem[16'h93C6] = 8'h48;
mem[16'h93C7] = 8'h00;
mem[16'h93C8] = 8'h00;
mem[16'h93C9] = 8'h0C;
mem[16'h93CA] = 8'h60;
mem[16'h93CB] = 8'h00;
mem[16'h93CC] = 8'h00;
mem[16'h93CD] = 8'h71;
mem[16'h93CE] = 8'h00;
mem[16'h93CF] = 8'h03;
mem[16'h93D0] = 8'h00;
mem[16'h93D1] = 8'h71;
mem[16'h93D2] = 8'h00;
mem[16'h93D3] = 8'h03;
mem[16'h93D4] = 8'h00;
mem[16'h93D5] = 8'h71;
mem[16'h93D6] = 8'h00;
mem[16'h93D7] = 8'h03;
mem[16'h93D8] = 8'h00;
mem[16'h93D9] = 8'h0C;
mem[16'h93DA] = 8'h60;
mem[16'h93DB] = 8'h00;
mem[16'h93DC] = 8'h00;
mem[16'h93DD] = 8'h60;
mem[16'h93DE] = 8'h48;
mem[16'h93DF] = 8'h00;
mem[16'h93E0] = 8'h00;
mem[16'h93E1] = 8'h20;
mem[16'h93E2] = 8'h11;
mem[16'h93E3] = 8'h00;
mem[16'h93E4] = 8'h00;
mem[16'h93E5] = 8'h20;
mem[16'h93E6] = 8'h00;
mem[16'h93E7] = 8'h00;
mem[16'h93E8] = 8'h00;
mem[16'h93E9] = 8'h00;
mem[16'h93EA] = 8'h22;
mem[16'h93EB] = 8'h00;
mem[16'h93EC] = 8'h00;
mem[16'h93ED] = 8'h00;
mem[16'h93EE] = 8'h16;
mem[16'h93EF] = 8'h01;
mem[16'h93F0] = 8'h00;
mem[16'h93F1] = 8'h40;
mem[16'h93F2] = 8'h00;
mem[16'h93F3] = 8'h01;
mem[16'h93F4] = 8'h00;
mem[16'h93F5] = 8'h40;
mem[16'h93F6] = 8'h00;
mem[16'h93F7] = 8'h04;
mem[16'h93F8] = 8'h00;
mem[16'h93F9] = 8'h00;
mem[16'h93FA] = 8'h02;
mem[16'h93FB] = 8'h04;
mem[16'h93FC] = 8'h00;
mem[16'h93FD] = 8'h00;
mem[16'h93FE] = 8'h08;
mem[16'h93FF] = 8'h04;
mem[16'h9400] = 8'h00;
mem[16'h9401] = 8'h00;
mem[16'h9402] = 8'h08;
mem[16'h9403] = 8'h10;
mem[16'h9404] = 8'h00;
mem[16'h9405] = 8'h00;
mem[16'h9406] = 8'h08;
mem[16'h9407] = 8'h40;
mem[16'h9408] = 8'h00;
mem[16'h9409] = 8'h00;
mem[16'h940A] = 8'h08;
mem[16'h940B] = 8'h00;
mem[16'h940C] = 8'h02;
mem[16'h940D] = 8'h00;
mem[16'h940E] = 8'h11;
mem[16'h940F] = 8'h00;
mem[16'h9410] = 8'h00;
mem[16'h9411] = 8'h00;
mem[16'h9412] = 8'h4B;
mem[16'h9413] = 8'h00;
mem[16'h9414] = 8'h00;
mem[16'h9415] = 8'h20;
mem[16'h9416] = 8'h40;
mem[16'h9417] = 8'h00;
mem[16'h9418] = 8'h00;
mem[16'h9419] = 8'h20;
mem[16'h941A] = 8'h00;
mem[16'h941B] = 8'h02;
mem[16'h941C] = 8'h00;
mem[16'h941D] = 8'h00;
mem[16'h941E] = 8'h01;
mem[16'h941F] = 8'h02;
mem[16'h9420] = 8'h00;
mem[16'h9421] = 8'h00;
mem[16'h9422] = 8'h04;
mem[16'h9423] = 8'h02;
mem[16'h9424] = 8'h00;
mem[16'h9425] = 8'h00;
mem[16'h9426] = 8'h04;
mem[16'h9427] = 8'h08;
mem[16'h9428] = 8'h00;
mem[16'h9429] = 8'h00;
mem[16'h942A] = 8'h04;
mem[16'h942B] = 8'h20;
mem[16'h942C] = 8'h00;
mem[16'h942D] = 8'h00;
mem[16'h942E] = 8'h04;
mem[16'h942F] = 8'h00;
mem[16'h9430] = 8'h01;
mem[16'h9431] = 8'h40;
mem[16'h9432] = 8'h08;
mem[16'h9433] = 8'h00;
mem[16'h9434] = 8'h00;
mem[16'h9435] = 8'h40;
mem[16'h9436] = 8'h25;
mem[16'h9437] = 8'h00;
mem[16'h9438] = 8'h00;
mem[16'h9439] = 8'h10;
mem[16'h943A] = 8'h20;
mem[16'h943B] = 8'h00;
mem[16'h943C] = 8'h00;
mem[16'h943D] = 8'h10;
mem[16'h943E] = 8'h00;
mem[16'h943F] = 8'h01;
mem[16'h9440] = 8'h00;
mem[16'h9441] = 8'h40;
mem[16'h9442] = 8'h00;
mem[16'h9443] = 8'h01;
mem[16'h9444] = 8'h00;
mem[16'h9445] = 8'h00;
mem[16'h9446] = 8'h02;
mem[16'h9447] = 8'h01;
mem[16'h9448] = 8'h00;
mem[16'h9449] = 8'h00;
mem[16'h944A] = 8'h02;
mem[16'h944B] = 8'h04;
mem[16'h944C] = 8'h00;
mem[16'h944D] = 8'h00;
mem[16'h944E] = 8'h02;
mem[16'h944F] = 8'h10;
mem[16'h9450] = 8'h00;
mem[16'h9451] = 8'h00;
mem[16'h9452] = 8'h02;
mem[16'h9453] = 8'h40;
mem[16'h9454] = 8'h00;
mem[16'h9455] = 8'h20;
mem[16'h9456] = 8'h04;
mem[16'h9457] = 8'h00;
mem[16'h9458] = 8'h00;
mem[16'h9459] = 8'h60;
mem[16'h945A] = 8'h12;
mem[16'h945B] = 8'h00;
mem[16'h945C] = 8'h00;
mem[16'h945D] = 8'h08;
mem[16'h945E] = 8'h10;
mem[16'h945F] = 8'h00;
mem[16'h9460] = 8'h00;
mem[16'h9461] = 8'h08;
mem[16'h9462] = 8'h40;
mem[16'h9463] = 8'h00;
mem[16'h9464] = 8'h00;
mem[16'h9465] = 8'h20;
mem[16'h9466] = 8'h40;
mem[16'h9467] = 8'h00;
mem[16'h9468] = 8'h00;
mem[16'h9469] = 8'h00;
mem[16'h946A] = 8'h41;
mem[16'h946B] = 8'h00;
mem[16'h946C] = 8'h00;
mem[16'h946D] = 8'h00;
mem[16'h946E] = 8'h01;
mem[16'h946F] = 8'h02;
mem[16'h9470] = 8'h00;
mem[16'h9471] = 8'h00;
mem[16'h9472] = 8'h01;
mem[16'h9473] = 8'h08;
mem[16'h9474] = 8'h00;
mem[16'h9475] = 8'h00;
mem[16'h9476] = 8'h01;
mem[16'h9477] = 8'h20;
mem[16'h9478] = 8'h00;
mem[16'h9479] = 8'h10;
mem[16'h947A] = 8'h02;
mem[16'h947B] = 8'h00;
mem[16'h947C] = 8'h00;
mem[16'h947D] = 8'h30;
mem[16'h947E] = 8'h09;
mem[16'h947F] = 8'h00;
mem[16'h9480] = 8'h00;
mem[16'h9481] = 8'h04;
mem[16'h9482] = 8'h08;
mem[16'h9483] = 8'h00;
mem[16'h9484] = 8'h00;
mem[16'h9485] = 8'h04;
mem[16'h9486] = 8'h20;
mem[16'h9487] = 8'h00;
mem[16'h9488] = 8'h00;
mem[16'h9489] = 8'h10;
mem[16'h948A] = 8'h20;
mem[16'h948B] = 8'h00;
mem[16'h948C] = 8'h00;
mem[16'h948D] = 8'h40;
mem[16'h948E] = 8'h20;
mem[16'h948F] = 8'h00;
mem[16'h9490] = 8'h00;
mem[16'h9491] = 8'h40;
mem[16'h9492] = 8'h00;
mem[16'h9493] = 8'h01;
mem[16'h9494] = 8'h00;
mem[16'h9495] = 8'h40;
mem[16'h9496] = 8'h00;
mem[16'h9497] = 8'h04;
mem[16'h9498] = 8'h00;
mem[16'h9499] = 8'h40;
mem[16'h949A] = 8'h00;
mem[16'h949B] = 8'h10;
mem[16'h949C] = 8'h00;
mem[16'h949D] = 8'h08;
mem[16'h949E] = 8'h01;
mem[16'h949F] = 8'h00;
mem[16'h94A0] = 8'h00;
mem[16'h94A1] = 8'h58;
mem[16'h94A2] = 8'h04;
mem[16'h94A3] = 8'h00;
mem[16'h94A4] = 8'h00;
mem[16'h94A5] = 8'h02;
mem[16'h94A6] = 8'h04;
mem[16'h94A7] = 8'h00;
mem[16'h94A8] = 8'h00;
mem[16'h94A9] = 8'h02;
mem[16'h94AA] = 8'h10;
mem[16'h94AB] = 8'h00;
mem[16'h94AC] = 8'h00;
mem[16'h94AD] = 8'h08;
mem[16'h94AE] = 8'h10;
mem[16'h94AF] = 8'h00;
mem[16'h94B0] = 8'h00;
mem[16'h94B1] = 8'h20;
mem[16'h94B2] = 8'h10;
mem[16'h94B3] = 8'h00;
mem[16'h94B4] = 8'h00;
mem[16'h94B5] = 8'h20;
mem[16'h94B6] = 8'h40;
mem[16'h94B7] = 8'h00;
mem[16'h94B8] = 8'h00;
mem[16'h94B9] = 8'h20;
mem[16'h94BA] = 8'h00;
mem[16'h94BB] = 8'h02;
mem[16'h94BC] = 8'h00;
mem[16'h94BD] = 8'h20;
mem[16'h94BE] = 8'h00;
mem[16'h94BF] = 8'h08;
mem[16'h94C0] = 8'h00;
mem[16'h94C1] = 8'h44;
mem[16'h94C2] = 8'h00;
mem[16'h94C3] = 8'h00;
mem[16'h94C4] = 8'h00;
mem[16'h94C5] = 8'h2C;
mem[16'h94C6] = 8'h02;
mem[16'h94C7] = 8'h00;
mem[16'h94C8] = 8'h00;
mem[16'h94C9] = 8'h01;
mem[16'h94CA] = 8'h02;
mem[16'h94CB] = 8'h00;
mem[16'h94CC] = 8'h00;
mem[16'h94CD] = 8'h01;
mem[16'h94CE] = 8'h08;
mem[16'h94CF] = 8'h00;
mem[16'h94D0] = 8'h00;
mem[16'h94D1] = 8'h04;
mem[16'h94D2] = 8'h08;
mem[16'h94D3] = 8'h00;
mem[16'h94D4] = 8'h00;
mem[16'h94D5] = 8'h10;
mem[16'h94D6] = 8'h08;
mem[16'h94D7] = 8'h00;
mem[16'h94D8] = 8'h00;
mem[16'h94D9] = 8'h10;
mem[16'h94DA] = 8'h20;
mem[16'h94DB] = 8'h00;
mem[16'h94DC] = 8'h00;
mem[16'h94DD] = 8'h10;
mem[16'h94DE] = 8'h00;
mem[16'h94DF] = 8'h01;
mem[16'h94E0] = 8'h00;
mem[16'h94E1] = 8'h10;
mem[16'h94E2] = 8'h00;
mem[16'h94E3] = 8'h04;
mem[16'h94E4] = 8'h00;
mem[16'h94E5] = 8'h00;
mem[16'h94E6] = 8'h00;
mem[16'h94E7] = 8'h44;
mem[16'h94E8] = 8'h00;
mem[16'h94E9] = 8'h00;
mem[16'h94EA] = 8'h00;
mem[16'h94EB] = 8'h69;
mem[16'h94EC] = 8'h00;
mem[16'h94ED] = 8'h00;
mem[16'h94EE] = 8'h00;
mem[16'h94EF] = 8'h01;
mem[16'h94F0] = 8'h02;
mem[16'h94F1] = 8'h00;
mem[16'h94F2] = 8'h20;
mem[16'h94F3] = 8'h00;
mem[16'h94F4] = 8'h02;
mem[16'h94F5] = 8'h00;
mem[16'h94F6] = 8'h20;
mem[16'h94F7] = 8'h40;
mem[16'h94F8] = 8'h00;
mem[16'h94F9] = 8'h00;
mem[16'h94FA] = 8'h20;
mem[16'h94FB] = 8'h10;
mem[16'h94FC] = 8'h00;
mem[16'h94FD] = 8'h00;
mem[16'h94FE] = 8'h08;
mem[16'h94FF] = 8'h10;
mem[16'h9500] = 8'h00;
mem[16'h9501] = 8'h00;
mem[16'h9502] = 8'h02;
mem[16'h9503] = 8'h10;
mem[16'h9504] = 8'h00;
mem[16'h9505] = 8'h40;
mem[16'h9506] = 8'h00;
mem[16'h9507] = 8'h10;
mem[16'h9508] = 8'h00;
mem[16'h9509] = 8'h00;
mem[16'h950A] = 8'h00;
mem[16'h950B] = 8'h22;
mem[16'h950C] = 8'h00;
mem[16'h950D] = 8'h00;
mem[16'h950E] = 8'h40;
mem[16'h950F] = 8'h34;
mem[16'h9510] = 8'h00;
mem[16'h9511] = 8'h00;
mem[16'h9512] = 8'h40;
mem[16'h9513] = 8'h00;
mem[16'h9514] = 8'h01;
mem[16'h9515] = 8'h00;
mem[16'h9516] = 8'h10;
mem[16'h9517] = 8'h00;
mem[16'h9518] = 8'h01;
mem[16'h9519] = 8'h00;
mem[16'h951A] = 8'h10;
mem[16'h951B] = 8'h20;
mem[16'h951C] = 8'h00;
mem[16'h951D] = 8'h00;
mem[16'h951E] = 8'h10;
mem[16'h951F] = 8'h08;
mem[16'h9520] = 8'h00;
mem[16'h9521] = 8'h00;
mem[16'h9522] = 8'h04;
mem[16'h9523] = 8'h08;
mem[16'h9524] = 8'h00;
mem[16'h9525] = 8'h00;
mem[16'h9526] = 8'h01;
mem[16'h9527] = 8'h08;
mem[16'h9528] = 8'h00;
mem[16'h9529] = 8'h20;
mem[16'h952A] = 8'h00;
mem[16'h952B] = 8'h08;
mem[16'h952C] = 8'h00;
mem[16'h952D] = 8'h00;
mem[16'h952E] = 8'h00;
mem[16'h952F] = 8'h11;
mem[16'h9530] = 8'h00;
mem[16'h9531] = 8'h00;
mem[16'h9532] = 8'h20;
mem[16'h9533] = 8'h1A;
mem[16'h9534] = 8'h00;
mem[16'h9535] = 8'h00;
mem[16'h9536] = 8'h20;
mem[16'h9537] = 8'h40;
mem[16'h9538] = 8'h00;
mem[16'h9539] = 8'h00;
mem[16'h953A] = 8'h08;
mem[16'h953B] = 8'h40;
mem[16'h953C] = 8'h00;
mem[16'h953D] = 8'h00;
mem[16'h953E] = 8'h08;
mem[16'h953F] = 8'h10;
mem[16'h9540] = 8'h00;
mem[16'h9541] = 8'h00;
mem[16'h9542] = 8'h08;
mem[16'h9543] = 8'h04;
mem[16'h9544] = 8'h00;
mem[16'h9545] = 8'h00;
mem[16'h9546] = 8'h02;
mem[16'h9547] = 8'h04;
mem[16'h9548] = 8'h00;
mem[16'h9549] = 8'h40;
mem[16'h954A] = 8'h00;
mem[16'h954B] = 8'h04;
mem[16'h954C] = 8'h00;
mem[16'h954D] = 8'h10;
mem[16'h954E] = 8'h00;
mem[16'h954F] = 8'h04;
mem[16'h9550] = 8'h00;
mem[16'h9551] = 8'h00;
mem[16'h9552] = 8'h40;
mem[16'h9553] = 8'h08;
mem[16'h9554] = 8'h00;
mem[16'h9555] = 8'h00;
mem[16'h9556] = 8'h10;
mem[16'h9557] = 8'h0D;
mem[16'h9558] = 8'h00;
mem[16'h9559] = 8'h00;
mem[16'h955A] = 8'h10;
mem[16'h955B] = 8'h20;
mem[16'h955C] = 8'h00;
mem[16'h955D] = 8'h00;
mem[16'h955E] = 8'h04;
mem[16'h955F] = 8'h20;
mem[16'h9560] = 8'h00;
mem[16'h9561] = 8'h00;
mem[16'h9562] = 8'h04;
mem[16'h9563] = 8'h08;
mem[16'h9564] = 8'h00;
mem[16'h9565] = 8'h00;
mem[16'h9566] = 8'h04;
mem[16'h9567] = 8'h02;
mem[16'h9568] = 8'h00;
mem[16'h9569] = 8'h00;
mem[16'h956A] = 8'h01;
mem[16'h956B] = 8'h02;
mem[16'h956C] = 8'h00;
mem[16'h956D] = 8'h20;
mem[16'h956E] = 8'h00;
mem[16'h956F] = 8'h02;
mem[16'h9570] = 8'h00;
mem[16'h9571] = 8'h08;
mem[16'h9572] = 8'h00;
mem[16'h9573] = 8'h02;
mem[16'h9574] = 8'h00;
mem[16'h9575] = 8'h00;
mem[16'h9576] = 8'h20;
mem[16'h9577] = 8'h04;
mem[16'h9578] = 8'h00;
mem[16'h9579] = 8'h00;
mem[16'h957A] = 8'h48;
mem[16'h957B] = 8'h06;
mem[16'h957C] = 8'h00;
mem[16'h957D] = 8'h00;
mem[16'h957E] = 8'h08;
mem[16'h957F] = 8'h10;
mem[16'h9580] = 8'h00;
mem[16'h9581] = 8'h00;
mem[16'h9582] = 8'h02;
mem[16'h9583] = 8'h10;
mem[16'h9584] = 8'h00;
mem[16'h9585] = 8'h00;
mem[16'h9586] = 8'h02;
mem[16'h9587] = 8'h04;
mem[16'h9588] = 8'h00;
mem[16'h9589] = 8'h00;
mem[16'h958A] = 8'h02;
mem[16'h958B] = 8'h01;
mem[16'h958C] = 8'h00;
mem[16'h958D] = 8'h40;
mem[16'h958E] = 8'h00;
mem[16'h958F] = 8'h01;
mem[16'h9590] = 8'h00;
mem[16'h9591] = 8'h10;
mem[16'h9592] = 8'h00;
mem[16'h9593] = 8'h01;
mem[16'h9594] = 8'h00;
mem[16'h9595] = 8'h04;
mem[16'h9596] = 8'h00;
mem[16'h9597] = 8'h01;
mem[16'h9598] = 8'h00;
mem[16'h9599] = 8'h00;
mem[16'h959A] = 8'h10;
mem[16'h959B] = 8'h02;
mem[16'h959C] = 8'h00;
mem[16'h959D] = 8'h00;
mem[16'h959E] = 8'h24;
mem[16'h959F] = 8'h03;
mem[16'h95A0] = 8'h00;
mem[16'h95A1] = 8'h00;
mem[16'h95A2] = 8'h04;
mem[16'h95A3] = 8'h08;
mem[16'h95A4] = 8'h00;
mem[16'h95A5] = 8'h00;
mem[16'h95A6] = 8'h01;
mem[16'h95A7] = 8'h08;
mem[16'h95A8] = 8'h00;
mem[16'h95A9] = 8'h00;
mem[16'h95AA] = 8'h01;
mem[16'h95AB] = 8'h02;
mem[16'h95AC] = 8'h00;
mem[16'h95AD] = 8'h00;
mem[16'h95AE] = 8'h41;
mem[16'h95AF] = 8'h00;
mem[16'h95B0] = 8'h00;
mem[16'h95B1] = 8'h20;
mem[16'h95B2] = 8'h40;
mem[16'h95B3] = 8'h00;
mem[16'h95B4] = 8'h00;
mem[16'h95B5] = 8'h08;
mem[16'h95B6] = 8'h40;
mem[16'h95B7] = 8'h00;
mem[16'h95B8] = 8'h00;
mem[16'h95B9] = 8'h02;
mem[16'h95BA] = 8'h40;
mem[16'h95BB] = 8'h00;
mem[16'h95BC] = 8'h00;
mem[16'h95BD] = 8'h00;
mem[16'h95BE] = 8'h08;
mem[16'h95BF] = 8'h01;
mem[16'h95C0] = 8'h00;
mem[16'h95C1] = 8'h00;
mem[16'h95C2] = 8'h52;
mem[16'h95C3] = 8'h01;
mem[16'h95C4] = 8'h00;
mem[16'h95C5] = 8'h00;
mem[16'h95C6] = 8'h02;
mem[16'h95C7] = 8'h04;
mem[16'h95C8] = 8'h00;
mem[16'h95C9] = 8'h40;
mem[16'h95CA] = 8'h00;
mem[16'h95CB] = 8'h04;
mem[16'h95CC] = 8'h00;
mem[16'h95CD] = 8'h40;
mem[16'h95CE] = 8'h00;
mem[16'h95CF] = 8'h01;
mem[16'h95D0] = 8'h00;
mem[16'h95D1] = 8'h40;
mem[16'h95D2] = 8'h20;
mem[16'h95D3] = 8'h00;
mem[16'h95D4] = 8'h00;
mem[16'h95D5] = 8'h10;
mem[16'h95D6] = 8'h20;
mem[16'h95D7] = 8'h00;
mem[16'h95D8] = 8'h00;
mem[16'h95D9] = 8'h04;
mem[16'h95DA] = 8'h20;
mem[16'h95DB] = 8'h00;
mem[16'h95DC] = 8'h00;
mem[16'h95DD] = 8'h01;
mem[16'h95DE] = 8'h20;
mem[16'h95DF] = 8'h00;
mem[16'h95E0] = 8'h00;
mem[16'h95E1] = 8'h0D;
mem[16'h95E2] = 8'h13;
mem[16'h95E3] = 8'hE4;
mem[16'h95E4] = 8'h20;
mem[16'h95E5] = 8'h36;
mem[16'h95E6] = 8'h38;
mem[16'h95E7] = 8'h34;
mem[16'h95E8] = 8'h31;
mem[16'h95E9] = 8'h30;
mem[16'h95EA] = 8'h42;
mem[16'h95EB] = 8'h30;
mem[16'h95EC] = 8'h30;
mem[16'h95ED] = 8'h32;
mem[16'h95EE] = 8'h38;
mem[16'h95EF] = 8'h36;
mem[16'h95F0] = 8'h33;
mem[16'h95F1] = 8'h30;
mem[16'h95F2] = 8'h41;
mem[16'h95F3] = 8'h30;
mem[16'h95F4] = 8'h30;
mem[16'h95F5] = 8'h0D;
mem[16'h95F6] = 8'h13;
mem[16'h95F7] = 8'hE4;
mem[16'h95F8] = 8'h20;
mem[16'h95F9] = 8'h30;
mem[16'h95FA] = 8'h30;
mem[16'h95FB] = 8'h30;
mem[16'h95FC] = 8'h30;
mem[16'h95FD] = 8'h30;
mem[16'h95FE] = 8'h30;
mem[16'h95FF] = 8'h30;
mem[16'h9600] = 8'h30;
mem[16'h9601] = 8'h30;
mem[16'h9602] = 8'h30;
mem[16'h9603] = 8'h30;
mem[16'h9604] = 8'h30;
mem[16'h9605] = 8'h30;
mem[16'h9606] = 8'h30;
mem[16'h9607] = 8'h30;
mem[16'h9608] = 8'h30;
mem[16'h9609] = 8'h30;
mem[16'h960A] = 8'h30;
mem[16'h960B] = 8'h30;
mem[16'h960C] = 8'h30;
mem[16'h960D] = 8'h30;
mem[16'h960E] = 8'h30;
mem[16'h960F] = 8'h30;
mem[16'h9610] = 8'h30;
mem[16'h9611] = 8'h30;
mem[16'h9612] = 8'h30;
mem[16'h9613] = 8'h30;
mem[16'h9614] = 8'h30;
mem[16'h9615] = 8'h30;
mem[16'h9616] = 8'h30;
mem[16'h9617] = 8'h30;
mem[16'h9618] = 8'h30;
mem[16'h9619] = 8'h30;
mem[16'h961A] = 8'h30;
mem[16'h961B] = 8'h30;
mem[16'h961C] = 8'h30;
mem[16'h961D] = 8'h30;
mem[16'h961E] = 8'h30;
mem[16'h961F] = 8'h30;
mem[16'h9620] = 8'h30;
mem[16'h9621] = 8'h30;
mem[16'h9622] = 8'h30;
mem[16'h9623] = 8'h30;
mem[16'h9624] = 8'h30;
mem[16'h9625] = 8'h30;
mem[16'h9626] = 8'h30;
mem[16'h9627] = 8'h30;
mem[16'h9628] = 8'h30;
mem[16'h9629] = 8'h30;
mem[16'h962A] = 8'h30;
mem[16'h962B] = 8'h30;
mem[16'h962C] = 8'h30;
mem[16'h962D] = 8'h30;
mem[16'h962E] = 8'h30;
mem[16'h962F] = 8'h30;
mem[16'h9630] = 8'h30;
mem[16'h9631] = 8'h30;
mem[16'h9632] = 8'h30;
mem[16'h9633] = 8'h30;
mem[16'h9634] = 8'h30;
mem[16'h9635] = 8'h30;
mem[16'h9636] = 8'h30;
mem[16'h9637] = 8'h30;
mem[16'h9638] = 8'h30;
mem[16'h9639] = 8'h30;
mem[16'h963A] = 8'h30;
mem[16'h963B] = 8'h30;
mem[16'h963C] = 8'h30;
mem[16'h963D] = 8'h30;
mem[16'h963E] = 8'h30;
mem[16'h963F] = 8'h30;
mem[16'h9640] = 8'h30;
mem[16'h9641] = 8'h30;
mem[16'h9642] = 8'h30;
mem[16'h9643] = 8'h30;
mem[16'h9644] = 8'h30;
mem[16'h9645] = 8'h30;
mem[16'h9646] = 8'h30;
mem[16'h9647] = 8'h30;
mem[16'h9648] = 8'h30;
mem[16'h9649] = 8'h30;
mem[16'h964A] = 8'h30;
mem[16'h964B] = 8'h30;
mem[16'h964C] = 8'h30;
mem[16'h964D] = 8'h30;
mem[16'h964E] = 8'h30;
mem[16'h964F] = 8'h30;
mem[16'h9650] = 8'h30;
mem[16'h9651] = 8'h30;
mem[16'h9652] = 8'h30;
mem[16'h9653] = 8'h30;
mem[16'h9654] = 8'h30;
mem[16'h9655] = 8'h30;
mem[16'h9656] = 8'h30;
mem[16'h9657] = 8'h30;
mem[16'h9658] = 8'h30;
mem[16'h9659] = 8'h30;
mem[16'h965A] = 8'h30;
mem[16'h965B] = 8'h30;
mem[16'h965C] = 8'h30;
mem[16'h965D] = 8'h30;
mem[16'h965E] = 8'h30;
mem[16'h965F] = 8'h30;
mem[16'h9660] = 8'h30;
mem[16'h9661] = 8'h30;
mem[16'h9662] = 8'h30;
mem[16'h9663] = 8'h30;
mem[16'h9664] = 8'h30;
mem[16'h9665] = 8'h30;
mem[16'h9666] = 8'h30;
mem[16'h9667] = 8'h30;
mem[16'h9668] = 8'h30;
mem[16'h9669] = 8'h30;
mem[16'h966A] = 8'h30;
mem[16'h966B] = 8'h30;
mem[16'h966C] = 8'h30;
mem[16'h966D] = 8'h30;
mem[16'h966E] = 8'h30;
mem[16'h966F] = 8'h30;
mem[16'h9670] = 8'h30;
mem[16'h9671] = 8'h30;
mem[16'h9672] = 8'h30;
mem[16'h9673] = 8'h30;
mem[16'h9674] = 8'h30;
mem[16'h9675] = 8'h30;
mem[16'h9676] = 8'h30;
mem[16'h9677] = 8'h30;
mem[16'h9678] = 8'h30;
mem[16'h9679] = 8'h30;
mem[16'h967A] = 8'h30;
mem[16'h967B] = 8'h30;
mem[16'h967C] = 8'h30;
mem[16'h967D] = 8'h30;
mem[16'h967E] = 8'h30;
mem[16'h967F] = 8'h30;
mem[16'h9680] = 8'h30;
mem[16'h9681] = 8'h30;
mem[16'h9682] = 8'h30;
mem[16'h9683] = 8'h30;
mem[16'h9684] = 8'h30;
mem[16'h9685] = 8'h30;
mem[16'h9686] = 8'h30;
mem[16'h9687] = 8'h30;
mem[16'h9688] = 8'h30;
mem[16'h9689] = 8'h30;
mem[16'h968A] = 8'h30;
mem[16'h968B] = 8'h30;
mem[16'h968C] = 8'h30;
mem[16'h968D] = 8'h30;
mem[16'h968E] = 8'h30;
mem[16'h968F] = 8'h30;
mem[16'h9690] = 8'h30;
mem[16'h9691] = 8'h30;
mem[16'h9692] = 8'h30;
mem[16'h9693] = 8'h30;
mem[16'h9694] = 8'h30;
mem[16'h9695] = 8'h30;
mem[16'h9696] = 8'h30;
mem[16'h9697] = 8'h30;
mem[16'h9698] = 8'h30;
mem[16'h9699] = 8'h30;
mem[16'h969A] = 8'h30;
mem[16'h969B] = 8'h30;
mem[16'h969C] = 8'h30;
mem[16'h969D] = 8'h30;
mem[16'h969E] = 8'h30;
mem[16'h969F] = 8'h30;
mem[16'h96A0] = 8'h30;
mem[16'h96A1] = 8'h30;
mem[16'h96A2] = 8'h30;
mem[16'h96A3] = 8'h30;
mem[16'h96A4] = 8'h30;
mem[16'h96A5] = 8'h30;
mem[16'h96A6] = 8'h30;
mem[16'h96A7] = 8'h30;
mem[16'h96A8] = 8'h30;
mem[16'h96A9] = 8'h30;
mem[16'h96AA] = 8'h30;
mem[16'h96AB] = 8'h30;
mem[16'h96AC] = 8'h30;
mem[16'h96AD] = 8'h30;
mem[16'h96AE] = 8'h30;
mem[16'h96AF] = 8'h30;
mem[16'h96B0] = 8'h30;
mem[16'h96B1] = 8'h30;
mem[16'h96B2] = 8'h30;
mem[16'h96B3] = 8'h30;
mem[16'h96B4] = 8'h30;
mem[16'h96B5] = 8'h30;
mem[16'h96B6] = 8'h30;
mem[16'h96B7] = 8'h30;
mem[16'h96B8] = 8'h30;
mem[16'h96B9] = 8'h30;
mem[16'h96BA] = 8'h30;
mem[16'h96BB] = 8'h30;
mem[16'h96BC] = 8'h30;
mem[16'h96BD] = 8'h30;
mem[16'h96BE] = 8'h30;
mem[16'h96BF] = 8'h30;
mem[16'h96C0] = 8'h30;
mem[16'h96C1] = 8'h30;
mem[16'h96C2] = 8'h30;
mem[16'h96C3] = 8'h30;
mem[16'h96C4] = 8'h30;
mem[16'h96C5] = 8'h30;
mem[16'h96C6] = 8'h30;
mem[16'h96C7] = 8'h30;
mem[16'h96C8] = 8'h30;
mem[16'h96C9] = 8'h30;
mem[16'h96CA] = 8'h30;
mem[16'h96CB] = 8'h30;
mem[16'h96CC] = 8'h30;
mem[16'h96CD] = 8'h30;
mem[16'h96CE] = 8'h30;
mem[16'h96CF] = 8'h30;
mem[16'h96D0] = 8'h30;
mem[16'h96D1] = 8'h30;
mem[16'h96D2] = 8'h30;
mem[16'h96D3] = 8'h30;
mem[16'h96D4] = 8'h30;
mem[16'h96D5] = 8'h30;
mem[16'h96D6] = 8'h30;
mem[16'h96D7] = 8'h30;
mem[16'h96D8] = 8'h30;
mem[16'h96D9] = 8'h30;
mem[16'h96DA] = 8'h30;
mem[16'h96DB] = 8'h30;
mem[16'h96DC] = 8'h30;
mem[16'h96DD] = 8'h30;
mem[16'h96DE] = 8'h30;
mem[16'h96DF] = 8'h30;
mem[16'h96E0] = 8'h30;
mem[16'h96E1] = 8'h30;
mem[16'h96E2] = 8'h30;
mem[16'h96E3] = 8'h30;
mem[16'h96E4] = 8'h30;
mem[16'h96E5] = 8'h30;
mem[16'h96E6] = 8'h30;
mem[16'h96E7] = 8'h30;
mem[16'h96E8] = 8'h30;
mem[16'h96E9] = 8'h30;
mem[16'h96EA] = 8'h30;
mem[16'h96EB] = 8'h30;
mem[16'h96EC] = 8'h30;
mem[16'h96ED] = 8'h30;
mem[16'h96EE] = 8'h30;
mem[16'h96EF] = 8'h30;
mem[16'h96F0] = 8'h30;
mem[16'h96F1] = 8'h30;
mem[16'h96F2] = 8'h30;
mem[16'h96F3] = 8'h30;
mem[16'h96F4] = 8'h30;
mem[16'h96F5] = 8'h30;
mem[16'h96F6] = 8'h30;
mem[16'h96F7] = 8'h30;
mem[16'h96F8] = 8'h30;
mem[16'h96F9] = 8'h30;
mem[16'h96FA] = 8'h30;
mem[16'h96FB] = 8'h30;
mem[16'h96FC] = 8'h30;
mem[16'h96FD] = 8'h00;
mem[16'h96FE] = 8'h00;
mem[16'h96FF] = 8'h00;
mem[16'h9700] = 8'hA0;
mem[16'h9701] = 8'h03;
mem[16'h9702] = 8'h84;
mem[16'h9703] = 8'h37;
mem[16'h9704] = 8'hA0;
mem[16'h9705] = 8'h09;
mem[16'h9706] = 8'h84;
mem[16'h9707] = 8'h36;
mem[16'h9708] = 8'h60;
mem[16'h9709] = 8'h48;
mem[16'h970A] = 8'h84;
mem[16'h970B] = 8'h4E;
mem[16'h970C] = 8'hC9;
mem[16'h970D] = 8'h8D;
mem[16'h970E] = 8'hF0;
mem[16'h970F] = 8'h68;
mem[16'h9710] = 8'hA5;
mem[16'h9711] = 8'h25;
mem[16'h9712] = 8'h4A;
mem[16'h9713] = 8'h29;
mem[16'h9714] = 8'h03;
mem[16'h9715] = 8'h09;
mem[16'h9716] = 8'h20;
mem[16'h9717] = 8'h85;
mem[16'h9718] = 8'h2B;
mem[16'h9719] = 8'hA5;
mem[16'h971A] = 8'h25;
mem[16'h971B] = 8'h6A;
mem[16'h971C] = 8'h08;
mem[16'h971D] = 8'h0A;
mem[16'h971E] = 8'h29;
mem[16'h971F] = 8'h18;
mem[16'h9720] = 8'h85;
mem[16'h9721] = 8'h2A;
mem[16'h9722] = 8'h0A;
mem[16'h9723] = 8'h0A;
mem[16'h9724] = 8'h05;
mem[16'h9725] = 8'h2A;
mem[16'h9726] = 8'h0A;
mem[16'h9727] = 8'h28;
mem[16'h9728] = 8'h6A;
mem[16'h9729] = 8'h18;
mem[16'h972A] = 8'h65;
mem[16'h972B] = 8'h24;
mem[16'h972C] = 8'h85;
mem[16'h972D] = 8'h2A;
mem[16'h972E] = 8'h68;
mem[16'h972F] = 8'h29;
mem[16'h9730] = 8'h7F;
mem[16'h9731] = 8'h48;
mem[16'h9732] = 8'hA9;
mem[16'h9733] = 8'h00;
mem[16'h9734] = 8'h85;
mem[16'h9735] = 8'h27;
mem[16'h9736] = 8'h68;
mem[16'h9737] = 8'h48;
mem[16'h9738] = 8'h2A;
mem[16'h9739] = 8'h26;
mem[16'h973A] = 8'h27;
mem[16'h973B] = 8'h2A;
mem[16'h973C] = 8'h26;
mem[16'h973D] = 8'h27;
mem[16'h973E] = 8'h2A;
mem[16'h973F] = 8'h26;
mem[16'h9740] = 8'h27;
mem[16'h9741] = 8'h85;
mem[16'h9742] = 8'h26;
mem[16'h9743] = 8'hA5;
mem[16'h9744] = 8'h27;
mem[16'h9745] = 8'h18;
mem[16'h9746] = 8'h69;
mem[16'h9747] = 8'h04;
mem[16'h9748] = 8'h85;
mem[16'h9749] = 8'h27;
mem[16'h974A] = 8'hA0;
mem[16'h974B] = 8'h00;
mem[16'h974C] = 8'hB1;
mem[16'h974D] = 8'h26;
mem[16'h974E] = 8'h48;
mem[16'h974F] = 8'h84;
mem[16'h9750] = 8'h4F;
mem[16'h9751] = 8'hA0;
mem[16'h9752] = 8'h00;
mem[16'h9753] = 8'h51;
mem[16'h9754] = 8'h2A;
mem[16'h9755] = 8'h91;
mem[16'h9756] = 8'h2A;
mem[16'h9757] = 8'hA5;
mem[16'h9758] = 8'h2B;
mem[16'h9759] = 8'hEA;
mem[16'h975A] = 8'hEA;
mem[16'h975B] = 8'h85;
mem[16'h975C] = 8'h2B;
mem[16'h975D] = 8'h68;
mem[16'h975E] = 8'h51;
mem[16'h975F] = 8'h2A;
mem[16'h9760] = 8'hEA;
mem[16'h9761] = 8'hEA;
mem[16'h9762] = 8'hA4;
mem[16'h9763] = 8'h4F;
mem[16'h9764] = 8'hA5;
mem[16'h9765] = 8'h2B;
mem[16'h9766] = 8'h18;
mem[16'h9767] = 8'h69;
mem[16'h9768] = 8'h04;
mem[16'h9769] = 8'h85;
mem[16'h976A] = 8'h2B;
mem[16'h976B] = 8'hC8;
mem[16'h976C] = 8'hC0;
mem[16'h976D] = 8'h08;
mem[16'h976E] = 8'hD0;
mem[16'h976F] = 8'hDC;
mem[16'h9770] = 8'hE6;
mem[16'h9771] = 8'h24;
mem[16'h9772] = 8'hA5;
mem[16'h9773] = 8'h24;
mem[16'h9774] = 8'hC5;
mem[16'h9775] = 8'h21;
mem[16'h9776] = 8'h90;
mem[16'h9777] = 8'h10;
mem[16'h9778] = 8'hA5;
mem[16'h9779] = 8'h20;
mem[16'h977A] = 8'h85;
mem[16'h977B] = 8'h24;
mem[16'h977C] = 8'hE6;
mem[16'h977D] = 8'h25;
mem[16'h977E] = 8'hA5;
mem[16'h977F] = 8'h25;
mem[16'h9780] = 8'hC5;
mem[16'h9781] = 8'h23;
mem[16'h9782] = 8'h90;
mem[16'h9783] = 8'h04;
mem[16'h9784] = 8'hA5;
mem[16'h9785] = 8'h22;
mem[16'h9786] = 8'h85;
mem[16'h9787] = 8'h25;
mem[16'h9788] = 8'hA4;
mem[16'h9789] = 8'h4E;
mem[16'h978A] = 8'h68;
mem[16'h978B] = 8'h60;
mem[16'h978C] = 8'hFF;
mem[16'h978D] = 8'hFF;
mem[16'h978E] = 8'h00;
mem[16'h978F] = 8'h00;
mem[16'h9790] = 8'hFF;
mem[16'h9791] = 8'hFF;
mem[16'h9792] = 8'h00;
mem[16'h9793] = 8'h00;
mem[16'h9794] = 8'hFF;
mem[16'h9795] = 8'hFF;
mem[16'h9796] = 8'h00;
mem[16'h9797] = 8'h00;
mem[16'h9798] = 8'hFF;
mem[16'h9799] = 8'hFF;
mem[16'h979A] = 8'h00;
mem[16'h979B] = 8'h00;
mem[16'h979C] = 8'hFF;
mem[16'h979D] = 8'hFF;
mem[16'h979E] = 8'h00;
mem[16'h979F] = 8'h00;
mem[16'h97A0] = 8'hFF;
mem[16'h97A1] = 8'hFF;
mem[16'h97A2] = 8'h00;
mem[16'h97A3] = 8'h00;
mem[16'h97A4] = 8'hFF;
mem[16'h97A5] = 8'hFF;
mem[16'h97A6] = 8'h00;
mem[16'h97A7] = 8'h00;
mem[16'h97A8] = 8'hFF;
mem[16'h97A9] = 8'hFF;
mem[16'h97AA] = 8'h00;
mem[16'h97AB] = 8'h00;
mem[16'h97AC] = 8'hFF;
mem[16'h97AD] = 8'hFF;
mem[16'h97AE] = 8'h00;
mem[16'h97AF] = 8'h00;
mem[16'h97B0] = 8'hFF;
mem[16'h97B1] = 8'hFF;
mem[16'h97B2] = 8'h00;
mem[16'h97B3] = 8'h00;
mem[16'h97B4] = 8'hFF;
mem[16'h97B5] = 8'hFF;
mem[16'h97B6] = 8'h00;
mem[16'h97B7] = 8'h00;
mem[16'h97B8] = 8'hFF;
mem[16'h97B9] = 8'hFF;
mem[16'h97BA] = 8'h00;
mem[16'h97BB] = 8'h00;
mem[16'h97BC] = 8'hFF;
mem[16'h97BD] = 8'hFF;
mem[16'h97BE] = 8'h00;
mem[16'h97BF] = 8'h00;
mem[16'h97C0] = 8'h00;
mem[16'h97C1] = 8'h00;
mem[16'h97C2] = 8'h00;
mem[16'h97C3] = 8'h00;
mem[16'h97C4] = 8'h00;
mem[16'h97C5] = 8'h00;
mem[16'h97C6] = 8'h00;
mem[16'h97C7] = 8'h00;
mem[16'h97C8] = 8'h00;
mem[16'h97C9] = 8'h00;
mem[16'h97CA] = 8'h00;
mem[16'h97CB] = 8'h00;
mem[16'h97CC] = 8'hB6;
mem[16'h97CD] = 8'h00;
mem[16'h97CE] = 8'h00;
mem[16'h97CF] = 8'h00;
mem[16'h97D0] = 8'h4C;
mem[16'h97D1] = 8'hBF;
mem[16'h97D2] = 8'h9D;
mem[16'h97D3] = 8'h4C;
mem[16'h97D4] = 8'h84;
mem[16'h97D5] = 8'h9D;
mem[16'h97D6] = 8'h4C;
mem[16'h97D7] = 8'hFD;
mem[16'h97D8] = 8'hAA;
mem[16'h97D9] = 8'h4C;
mem[16'h97DA] = 8'hB5;
mem[16'h97DB] = 8'hB7;
mem[16'h97DC] = 8'hAD;
mem[16'h97DD] = 8'h0F;
mem[16'h97DE] = 8'h9D;
mem[16'h97DF] = 8'hAC;
mem[16'h97E0] = 8'h0E;
mem[16'h97E1] = 8'h9D;
mem[16'h97E2] = 8'h60;
mem[16'h97E3] = 8'hAD;
mem[16'h97E4] = 8'hC2;
mem[16'h97E5] = 8'hAA;
mem[16'h97E6] = 8'hAC;
mem[16'h97E7] = 8'hC1;
mem[16'h97E8] = 8'hAA;
mem[16'h97E9] = 8'h60;
mem[16'h97EA] = 8'h4C;
mem[16'h97EB] = 8'h51;
mem[16'h97EC] = 8'hA8;
mem[16'h97ED] = 8'hEA;
mem[16'h97EE] = 8'hEA;
mem[16'h97EF] = 8'h4C;
mem[16'h97F0] = 8'h59;
mem[16'h97F1] = 8'hFA;
mem[16'h97F2] = 8'h43;
mem[16'h97F3] = 8'h30;
mem[16'h97F4] = 8'h95;
mem[16'h97F5] = 8'h4C;
mem[16'h97F6] = 8'h58;
mem[16'h97F7] = 8'hFF;
mem[16'h97F8] = 8'h4C;
mem[16'h97F9] = 8'h65;
mem[16'h97FA] = 8'hFF;
mem[16'h97FB] = 8'h4C;
mem[16'h97FC] = 8'h65;
mem[16'h97FD] = 8'hFF;
mem[16'h97FE] = 8'h65;
mem[16'h97FF] = 8'hFF;
mem[16'h9800] = 8'h00;
mem[16'h9801] = 8'hFF;
mem[16'h9802] = 8'hFF;
mem[16'h9803] = 8'h00;
mem[16'h9804] = 8'h00;
mem[16'h9805] = 8'hFF;
mem[16'h9806] = 8'hFF;
mem[16'h9807] = 8'h00;
mem[16'h9808] = 8'h00;
mem[16'h9809] = 8'hFF;
mem[16'h980A] = 8'hFF;
mem[16'h980B] = 8'h00;
mem[16'h980C] = 8'h00;
mem[16'h980D] = 8'hFF;
mem[16'h980E] = 8'hFF;
mem[16'h980F] = 8'h00;
mem[16'h9810] = 8'h00;
mem[16'h9811] = 8'hFF;
mem[16'h9812] = 8'hFF;
mem[16'h9813] = 8'h00;
mem[16'h9814] = 8'h00;
mem[16'h9815] = 8'hFF;
mem[16'h9816] = 8'hFF;
mem[16'h9817] = 8'h00;
mem[16'h9818] = 8'h00;
mem[16'h9819] = 8'hFF;
mem[16'h981A] = 8'hFF;
mem[16'h981B] = 8'h00;
mem[16'h981C] = 8'h00;
mem[16'h981D] = 8'hFF;
mem[16'h981E] = 8'hFF;
mem[16'h981F] = 8'h00;
mem[16'h9820] = 8'h00;
mem[16'h9821] = 8'hFF;
mem[16'h9822] = 8'hFF;
mem[16'h9823] = 8'h00;
mem[16'h9824] = 8'h00;
mem[16'h9825] = 8'hFF;
mem[16'h9826] = 8'hFF;
mem[16'h9827] = 8'h00;
mem[16'h9828] = 8'h00;
mem[16'h9829] = 8'hFF;
mem[16'h982A] = 8'hFF;
mem[16'h982B] = 8'h00;
mem[16'h982C] = 8'h00;
mem[16'h982D] = 8'hFF;
mem[16'h982E] = 8'hFF;
mem[16'h982F] = 8'h00;
mem[16'h9830] = 8'h00;
mem[16'h9831] = 8'hFF;
mem[16'h9832] = 8'hFF;
mem[16'h9833] = 8'h00;
mem[16'h9834] = 8'h00;
mem[16'h9835] = 8'hFF;
mem[16'h9836] = 8'hFF;
mem[16'h9837] = 8'h00;
mem[16'h9838] = 8'h00;
mem[16'h9839] = 8'h14;
mem[16'h983A] = 8'h22;
mem[16'h983B] = 8'h22;
mem[16'h983C] = 8'h22;
mem[16'h983D] = 8'h41;
mem[16'h983E] = 8'h7F;
mem[16'h983F] = 8'h08;
mem[16'h9840] = 8'h10;
mem[16'h9841] = 8'h08;
mem[16'h9842] = 8'h04;
mem[16'h9843] = 8'h7E;
mem[16'h9844] = 8'h04;
mem[16'h9845] = 8'h08;
mem[16'h9846] = 8'h10;
mem[16'h9847] = 8'h00;
mem[16'h9848] = 8'h08;
mem[16'h9849] = 8'h10;
mem[16'h984A] = 8'h20;
mem[16'h984B] = 8'h7E;
mem[16'h984C] = 8'h20;
mem[16'h984D] = 8'h10;
mem[16'h984E] = 8'h08;
mem[16'h984F] = 8'h00;
mem[16'h9850] = 8'h08;
mem[16'h9851] = 8'h08;
mem[16'h9852] = 8'h08;
mem[16'h9853] = 8'h49;
mem[16'h9854] = 8'h2A;
mem[16'h9855] = 8'h1C;
mem[16'h9856] = 8'h08;
mem[16'h9857] = 8'h00;
mem[16'h9858] = 8'h08;
mem[16'h9859] = 8'h1C;
mem[16'h985A] = 8'h2A;
mem[16'h985B] = 8'h49;
mem[16'h985C] = 8'h08;
mem[16'h985D] = 8'h08;
mem[16'h985E] = 8'h08;
mem[16'h985F] = 8'h00;
mem[16'h9860] = 8'h08;
mem[16'h9861] = 8'h49;
mem[16'h9862] = 8'h2A;
mem[16'h9863] = 8'h1C;
mem[16'h9864] = 8'h49;
mem[16'h9865] = 8'h2A;
mem[16'h9866] = 8'h1C;
mem[16'h9867] = 8'h08;
mem[16'h9868] = 8'h40;
mem[16'h9869] = 8'h60;
mem[16'h986A] = 8'h70;
mem[16'h986B] = 8'h78;
mem[16'h986C] = 8'h70;
mem[16'h986D] = 8'h60;
mem[16'h986E] = 8'h40;
mem[16'h986F] = 8'h00;
mem[16'h9870] = 8'h40;
mem[16'h9871] = 8'h40;
mem[16'h9872] = 8'h20;
mem[16'h9873] = 8'h20;
mem[16'h9874] = 8'h13;
mem[16'h9875] = 8'h14;
mem[16'h9876] = 8'h0C;
mem[16'h9877] = 8'h08;
mem[16'h9878] = 8'h1A;
mem[16'h9879] = 8'h00;
mem[16'h987A] = 8'h00;
mem[16'h987B] = 8'h7C;
mem[16'h987C] = 8'h2A;
mem[16'h987D] = 8'h28;
mem[16'h987E] = 8'h34;
mem[16'h987F] = 8'h00;
mem[16'h9880] = 8'h36;
mem[16'h9881] = 8'h7F;
mem[16'h9882] = 8'h7F;
mem[16'h9883] = 8'h7F;
mem[16'h9884] = 8'h3E;
mem[16'h9885] = 8'h1C;
mem[16'h9886] = 8'h08;
mem[16'h9887] = 8'h00;
mem[16'h9888] = 8'h08;
mem[16'h9889] = 8'h1C;
mem[16'h988A] = 8'h3E;
mem[16'h988B] = 8'h7F;
mem[16'h988C] = 8'h3E;
mem[16'h988D] = 8'h1C;
mem[16'h988E] = 8'h08;
mem[16'h988F] = 8'h00;
mem[16'h9890] = 8'h08;
mem[16'h9891] = 8'h1C;
mem[16'h9892] = 8'h3E;
mem[16'h9893] = 8'h7F;
mem[16'h9894] = 8'h7F;
mem[16'h9895] = 8'h2A;
mem[16'h9896] = 8'h08;
mem[16'h9897] = 8'h00;
mem[16'h9898] = 8'h08;
mem[16'h9899] = 8'h1C;
mem[16'h989A] = 8'h1C;
mem[16'h989B] = 8'h2A;
mem[16'h989C] = 8'h7F;
mem[16'h989D] = 8'h7F;
mem[16'h989E] = 8'h2A;
mem[16'h989F] = 8'h08;
mem[16'h98A0] = 8'h3E;
mem[16'h98A1] = 8'h08;
mem[16'h98A2] = 8'h08;
mem[16'h98A3] = 8'h22;
mem[16'h98A4] = 8'h36;
mem[16'h98A5] = 8'h2A;
mem[16'h98A6] = 8'h22;
mem[16'h98A7] = 8'h00;
mem[16'h98A8] = 8'h00;
mem[16'h98A9] = 8'h22;
mem[16'h98AA] = 8'h14;
mem[16'h98AB] = 8'h08;
mem[16'h98AC] = 8'h14;
mem[16'h98AD] = 8'h22;
mem[16'h98AE] = 8'h00;
mem[16'h98AF] = 8'h00;
mem[16'h98B0] = 8'h04;
mem[16'h98B1] = 8'h0E;
mem[16'h98B2] = 8'h04;
mem[16'h98B3] = 8'h04;
mem[16'h98B4] = 8'h00;
mem[16'h98B5] = 8'h00;
mem[16'h98B6] = 8'h00;
mem[16'h98B7] = 8'h00;
mem[16'h98B8] = 8'h00;
mem[16'h98B9] = 8'h08;
mem[16'h98BA] = 8'h00;
mem[16'h98BB] = 8'h3E;
mem[16'h98BC] = 8'h00;
mem[16'h98BD] = 8'h08;
mem[16'h98BE] = 8'h00;
mem[16'h98BF] = 8'h00;
mem[16'h98C0] = 8'h18;
mem[16'h98C1] = 8'h24;
mem[16'h98C2] = 8'h08;
mem[16'h98C3] = 8'h14;
mem[16'h98C4] = 8'h08;
mem[16'h98C5] = 8'h12;
mem[16'h98C6] = 8'h0C;
mem[16'h98C7] = 8'h00;
mem[16'h98C8] = 8'h10;
mem[16'h98C9] = 8'h38;
mem[16'h98CA] = 8'h04;
mem[16'h98CB] = 8'h04;
mem[16'h98CC] = 8'h38;
mem[16'h98CD] = 8'h10;
mem[16'h98CE] = 8'h00;
mem[16'h98CF] = 8'h00;
mem[16'h98D0] = 8'h08;
mem[16'h98D1] = 8'h1C;
mem[16'h98D2] = 8'h08;
mem[16'h98D3] = 8'h1C;
mem[16'h98D4] = 8'h3E;
mem[16'h98D5] = 8'h1C;
mem[16'h98D6] = 8'h3E;
mem[16'h98D7] = 8'h7F;
mem[16'h98D8] = 8'h08;
mem[16'h98D9] = 8'h3E;
mem[16'h98DA] = 8'h1C;
mem[16'h98DB] = 8'h08;
mem[16'h98DC] = 8'h1C;
mem[16'h98DD] = 8'h1C;
mem[16'h98DE] = 8'h3E;
mem[16'h98DF] = 8'h7F;
mem[16'h98E0] = 8'h00;
mem[16'h98E1] = 8'h2A;
mem[16'h98E2] = 8'h3E;
mem[16'h98E3] = 8'h1C;
mem[16'h98E4] = 8'h1C;
mem[16'h98E5] = 8'h1C;
mem[16'h98E6] = 8'h3E;
mem[16'h98E7] = 8'h7F;
mem[16'h98E8] = 8'h00;
mem[16'h98E9] = 8'h10;
mem[16'h98EA] = 8'h3C;
mem[16'h98EB] = 8'h3E;
mem[16'h98EC] = 8'h18;
mem[16'h98ED] = 8'h0C;
mem[16'h98EE] = 8'h1E;
mem[16'h98EF] = 8'h3F;
mem[16'h98F0] = 8'h00;
mem[16'h98F1] = 8'h08;
mem[16'h98F2] = 8'h18;
mem[16'h98F3] = 8'h3A;
mem[16'h98F4] = 8'h7B;
mem[16'h98F5] = 8'h3E;
mem[16'h98F6] = 8'h1C;
mem[16'h98F7] = 8'h7F;
mem[16'h98F8] = 8'h04;
mem[16'h98F9] = 8'h00;
mem[16'h98FA] = 8'h08;
mem[16'h98FB] = 8'h1C;
mem[16'h98FC] = 8'h1C;
mem[16'h98FD] = 8'h08;
mem[16'h98FE] = 8'h1C;
mem[16'h98FF] = 8'h3E;
mem[16'h9900] = 8'h00;
mem[16'h9901] = 8'h00;
mem[16'h9902] = 8'h00;
mem[16'h9903] = 8'h00;
mem[16'h9904] = 8'h00;
mem[16'h9905] = 8'h00;
mem[16'h9906] = 8'h00;
mem[16'h9907] = 8'h00;
mem[16'h9908] = 8'h10;
mem[16'h9909] = 8'h10;
mem[16'h990A] = 8'h10;
mem[16'h990B] = 8'h10;
mem[16'h990C] = 8'h00;
mem[16'h990D] = 8'h00;
mem[16'h990E] = 8'h10;
mem[16'h990F] = 8'h00;
mem[16'h9910] = 8'h24;
mem[16'h9911] = 8'h24;
mem[16'h9912] = 8'h24;
mem[16'h9913] = 8'h00;
mem[16'h9914] = 8'h00;
mem[16'h9915] = 8'h00;
mem[16'h9916] = 8'h00;
mem[16'h9917] = 8'h00;
mem[16'h9918] = 8'h24;
mem[16'h9919] = 8'h24;
mem[16'h991A] = 8'h7E;
mem[16'h991B] = 8'h24;
mem[16'h991C] = 8'h7E;
mem[16'h991D] = 8'h24;
mem[16'h991E] = 8'h24;
mem[16'h991F] = 8'h00;
mem[16'h9920] = 8'h10;
mem[16'h9921] = 8'h78;
mem[16'h9922] = 8'h14;
mem[16'h9923] = 8'h38;
mem[16'h9924] = 8'h50;
mem[16'h9925] = 8'h3C;
mem[16'h9926] = 8'h10;
mem[16'h9927] = 8'h00;
mem[16'h9928] = 8'h00;
mem[16'h9929] = 8'h46;
mem[16'h992A] = 8'h26;
mem[16'h992B] = 8'h10;
mem[16'h992C] = 8'h08;
mem[16'h992D] = 8'h64;
mem[16'h992E] = 8'h62;
mem[16'h992F] = 8'h00;
mem[16'h9930] = 8'h0C;
mem[16'h9931] = 8'h12;
mem[16'h9932] = 8'h12;
mem[16'h9933] = 8'h0C;
mem[16'h9934] = 8'h52;
mem[16'h9935] = 8'h22;
mem[16'h9936] = 8'h5C;
mem[16'h9937] = 8'h00;
mem[16'h9938] = 8'h20;
mem[16'h9939] = 8'h10;
mem[16'h993A] = 8'h08;
mem[16'h993B] = 8'h00;
mem[16'h993C] = 8'h00;
mem[16'h993D] = 8'h00;
mem[16'h993E] = 8'h00;
mem[16'h993F] = 8'h00;
mem[16'h9940] = 8'h20;
mem[16'h9941] = 8'h10;
mem[16'h9942] = 8'h08;
mem[16'h9943] = 8'h08;
mem[16'h9944] = 8'h08;
mem[16'h9945] = 8'h10;
mem[16'h9946] = 8'h20;
mem[16'h9947] = 8'h00;
mem[16'h9948] = 8'h04;
mem[16'h9949] = 8'h08;
mem[16'h994A] = 8'h10;
mem[16'h994B] = 8'h10;
mem[16'h994C] = 8'h10;
mem[16'h994D] = 8'h08;
mem[16'h994E] = 8'h04;
mem[16'h994F] = 8'h00;
mem[16'h9950] = 8'h10;
mem[16'h9951] = 8'h54;
mem[16'h9952] = 8'h38;
mem[16'h9953] = 8'h7C;
mem[16'h9954] = 8'h38;
mem[16'h9955] = 8'h54;
mem[16'h9956] = 8'h10;
mem[16'h9957] = 8'h00;
mem[16'h9958] = 8'h00;
mem[16'h9959] = 8'h10;
mem[16'h995A] = 8'h10;
mem[16'h995B] = 8'h7C;
mem[16'h995C] = 8'h10;
mem[16'h995D] = 8'h10;
mem[16'h995E] = 8'h00;
mem[16'h995F] = 8'h00;
mem[16'h9960] = 8'h00;
mem[16'h9961] = 8'h00;
mem[16'h9962] = 8'h00;
mem[16'h9963] = 8'h00;
mem[16'h9964] = 8'h00;
mem[16'h9965] = 8'h18;
mem[16'h9966] = 8'h18;
mem[16'h9967] = 8'h0C;
mem[16'h9968] = 8'h00;
mem[16'h9969] = 8'h00;
mem[16'h996A] = 8'h00;
mem[16'h996B] = 8'h7E;
mem[16'h996C] = 8'h00;
mem[16'h996D] = 8'h00;
mem[16'h996E] = 8'h00;
mem[16'h996F] = 8'h00;
mem[16'h9970] = 8'h00;
mem[16'h9971] = 8'h00;
mem[16'h9972] = 8'h00;
mem[16'h9973] = 8'h00;
mem[16'h9974] = 8'h00;
mem[16'h9975] = 8'h18;
mem[16'h9976] = 8'h18;
mem[16'h9977] = 8'h00;
mem[16'h9978] = 8'h28;
mem[16'h9979] = 8'h40;
mem[16'h997A] = 8'h20;
mem[16'h997B] = 8'h10;
mem[16'h997C] = 8'h08;
mem[16'h997D] = 8'h04;
mem[16'h997E] = 8'h02;
mem[16'h997F] = 8'h00;
mem[16'h9980] = 8'h3C;
mem[16'h9981] = 8'h42;
mem[16'h9982] = 8'h42;
mem[16'h9983] = 8'h42;
mem[16'h9984] = 8'h42;
mem[16'h9985] = 8'h42;
mem[16'h9986] = 8'h3C;
mem[16'h9987] = 8'h00;
mem[16'h9988] = 8'h10;
mem[16'h9989] = 8'h18;
mem[16'h998A] = 8'h14;
mem[16'h998B] = 8'h10;
mem[16'h998C] = 8'h10;
mem[16'h998D] = 8'h10;
mem[16'h998E] = 8'h7C;
mem[16'h998F] = 8'h00;
mem[16'h9990] = 8'h3C;
mem[16'h9991] = 8'h42;
mem[16'h9992] = 8'h40;
mem[16'h9993] = 8'h30;
mem[16'h9994] = 8'h0C;
mem[16'h9995] = 8'h02;
mem[16'h9996] = 8'h7E;
mem[16'h9997] = 8'h00;
mem[16'h9998] = 8'h3C;
mem[16'h9999] = 8'h42;
mem[16'h999A] = 8'h40;
mem[16'h999B] = 8'h38;
mem[16'h999C] = 8'h40;
mem[16'h999D] = 8'h42;
mem[16'h999E] = 8'h3C;
mem[16'h999F] = 8'h00;
mem[16'h99A0] = 8'h20;
mem[16'h99A1] = 8'h30;
mem[16'h99A2] = 8'h28;
mem[16'h99A3] = 8'h24;
mem[16'h99A4] = 8'h7E;
mem[16'h99A5] = 8'h20;
mem[16'h99A6] = 8'h20;
mem[16'h99A7] = 8'h00;
mem[16'h99A8] = 8'h7E;
mem[16'h99A9] = 8'h02;
mem[16'h99AA] = 8'h1E;
mem[16'h99AB] = 8'h20;
mem[16'h99AC] = 8'h40;
mem[16'h99AD] = 8'h22;
mem[16'h99AE] = 8'h1C;
mem[16'h99AF] = 8'h00;
mem[16'h99B0] = 8'h38;
mem[16'h99B1] = 8'h04;
mem[16'h99B2] = 8'h02;
mem[16'h99B3] = 8'h3E;
mem[16'h99B4] = 8'h42;
mem[16'h99B5] = 8'h42;
mem[16'h99B6] = 8'h3C;
mem[16'h99B7] = 8'h00;
mem[16'h99B8] = 8'h7E;
mem[16'h99B9] = 8'h42;
mem[16'h99BA] = 8'h20;
mem[16'h99BB] = 8'h10;
mem[16'h99BC] = 8'h08;
mem[16'h99BD] = 8'h08;
mem[16'h99BE] = 8'h08;
mem[16'h99BF] = 8'h00;
mem[16'h99C0] = 8'h3C;
mem[16'h99C1] = 8'h42;
mem[16'h99C2] = 8'h42;
mem[16'h99C3] = 8'h3C;
mem[16'h99C4] = 8'h42;
mem[16'h99C5] = 8'h42;
mem[16'h99C6] = 8'h3C;
mem[16'h99C7] = 8'h00;
mem[16'h99C8] = 8'h3C;
mem[16'h99C9] = 8'h42;
mem[16'h99CA] = 8'h42;
mem[16'h99CB] = 8'h7C;
mem[16'h99CC] = 8'h40;
mem[16'h99CD] = 8'h20;
mem[16'h99CE] = 8'h1C;
mem[16'h99CF] = 8'h00;
mem[16'h99D0] = 8'h00;
mem[16'h99D1] = 8'h00;
mem[16'h99D2] = 8'h18;
mem[16'h99D3] = 8'h18;
mem[16'h99D4] = 8'h00;
mem[16'h99D5] = 8'h18;
mem[16'h99D6] = 8'h18;
mem[16'h99D7] = 8'h00;
mem[16'h99D8] = 8'h00;
mem[16'h99D9] = 8'h00;
mem[16'h99DA] = 8'h18;
mem[16'h99DB] = 8'h18;
mem[16'h99DC] = 8'h00;
mem[16'h99DD] = 8'h18;
mem[16'h99DE] = 8'h18;
mem[16'h99DF] = 8'h0C;
mem[16'h99E0] = 8'h20;
mem[16'h99E1] = 8'h10;
mem[16'h99E2] = 8'h08;
mem[16'h99E3] = 8'h04;
mem[16'h99E4] = 8'h08;
mem[16'h99E5] = 8'h10;
mem[16'h99E6] = 8'h20;
mem[16'h99E7] = 8'h00;
mem[16'h99E8] = 8'h00;
mem[16'h99E9] = 8'h00;
mem[16'h99EA] = 8'h3E;
mem[16'h99EB] = 8'h00;
mem[16'h99EC] = 8'h3E;
mem[16'h99ED] = 8'h00;
mem[16'h99EE] = 8'h00;
mem[16'h99EF] = 8'h00;
mem[16'h99F0] = 8'h04;
mem[16'h99F1] = 8'h08;
mem[16'h99F2] = 8'h10;
mem[16'h99F3] = 8'h20;
mem[16'h99F4] = 8'h10;
mem[16'h99F5] = 8'h08;
mem[16'h99F6] = 8'h04;
mem[16'h99F7] = 8'h00;
mem[16'h99F8] = 8'h60;
mem[16'h99F9] = 8'h42;
mem[16'h99FA] = 8'h40;
mem[16'h99FB] = 8'h30;
mem[16'h99FC] = 8'h08;
mem[16'h99FD] = 8'h00;
mem[16'h99FE] = 8'h08;
mem[16'h99FF] = 8'h00;
mem[16'h9A00] = 8'h38;
mem[16'h9A01] = 8'h44;
mem[16'h9A02] = 8'h52;
mem[16'h9A03] = 8'h6A;
mem[16'h9A04] = 8'h32;
mem[16'h9A05] = 8'h04;
mem[16'h9A06] = 8'h78;
mem[16'h9A07] = 8'h00;
mem[16'h9A08] = 8'h18;
mem[16'h9A09] = 8'h24;
mem[16'h9A0A] = 8'h42;
mem[16'h9A0B] = 8'h7E;
mem[16'h9A0C] = 8'h42;
mem[16'h9A0D] = 8'h42;
mem[16'h9A0E] = 8'h42;
mem[16'h9A0F] = 8'h00;
mem[16'h9A10] = 8'h3E;
mem[16'h9A11] = 8'h44;
mem[16'h9A12] = 8'h44;
mem[16'h9A13] = 8'h3C;
mem[16'h9A14] = 8'h44;
mem[16'h9A15] = 8'h44;
mem[16'h9A16] = 8'h3E;
mem[16'h9A17] = 8'h00;
mem[16'h9A18] = 8'h3C;
mem[16'h9A19] = 8'h42;
mem[16'h9A1A] = 8'h02;
mem[16'h9A1B] = 8'h02;
mem[16'h9A1C] = 8'h02;
mem[16'h9A1D] = 8'h42;
mem[16'h9A1E] = 8'h3C;
mem[16'h9A1F] = 8'h00;
mem[16'h9A20] = 8'h3E;
mem[16'h9A21] = 8'h44;
mem[16'h9A22] = 8'h44;
mem[16'h9A23] = 8'h44;
mem[16'h9A24] = 8'h44;
mem[16'h9A25] = 8'h44;
mem[16'h9A26] = 8'h3E;
mem[16'h9A27] = 8'h00;
mem[16'h9A28] = 8'h7E;
mem[16'h9A29] = 8'h02;
mem[16'h9A2A] = 8'h02;
mem[16'h9A2B] = 8'h1E;
mem[16'h9A2C] = 8'h02;
mem[16'h9A2D] = 8'h02;
mem[16'h9A2E] = 8'h7E;
mem[16'h9A2F] = 8'h00;
mem[16'h9A30] = 8'h7E;
mem[16'h9A31] = 8'h02;
mem[16'h9A32] = 8'h02;
mem[16'h9A33] = 8'h1E;
mem[16'h9A34] = 8'h02;
mem[16'h9A35] = 8'h02;
mem[16'h9A36] = 8'h02;
mem[16'h9A37] = 8'h00;
mem[16'h9A38] = 8'h3C;
mem[16'h9A39] = 8'h42;
mem[16'h9A3A] = 8'h02;
mem[16'h9A3B] = 8'h72;
mem[16'h9A3C] = 8'h42;
mem[16'h9A3D] = 8'h42;
mem[16'h9A3E] = 8'h3C;
mem[16'h9A3F] = 8'h00;
mem[16'h9A40] = 8'h42;
mem[16'h9A41] = 8'h42;
mem[16'h9A42] = 8'h42;
mem[16'h9A43] = 8'h7E;
mem[16'h9A44] = 8'h42;
mem[16'h9A45] = 8'h42;
mem[16'h9A46] = 8'h42;
mem[16'h9A47] = 8'h00;
mem[16'h9A48] = 8'h38;
mem[16'h9A49] = 8'h10;
mem[16'h9A4A] = 8'h10;
mem[16'h9A4B] = 8'h10;
mem[16'h9A4C] = 8'h10;
mem[16'h9A4D] = 8'h10;
mem[16'h9A4E] = 8'h38;
mem[16'h9A4F] = 8'h00;
mem[16'h9A50] = 8'h70;
mem[16'h9A51] = 8'h20;
mem[16'h9A52] = 8'h20;
mem[16'h9A53] = 8'h20;
mem[16'h9A54] = 8'h20;
mem[16'h9A55] = 8'h22;
mem[16'h9A56] = 8'h1C;
mem[16'h9A57] = 8'h00;
mem[16'h9A58] = 8'h42;
mem[16'h9A59] = 8'h22;
mem[16'h9A5A] = 8'h12;
mem[16'h9A5B] = 8'h0E;
mem[16'h9A5C] = 8'h12;
mem[16'h9A5D] = 8'h22;
mem[16'h9A5E] = 8'h42;
mem[16'h9A5F] = 8'h00;
mem[16'h9A60] = 8'h02;
mem[16'h9A61] = 8'h02;
mem[16'h9A62] = 8'h02;
mem[16'h9A63] = 8'h02;
mem[16'h9A64] = 8'h02;
mem[16'h9A65] = 8'h02;
mem[16'h9A66] = 8'h7E;
mem[16'h9A67] = 8'h00;
mem[16'h9A68] = 8'h42;
mem[16'h9A69] = 8'h66;
mem[16'h9A6A] = 8'h5A;
mem[16'h9A6B] = 8'h5A;
mem[16'h9A6C] = 8'h42;
mem[16'h9A6D] = 8'h42;
mem[16'h9A6E] = 8'h42;
mem[16'h9A6F] = 8'h00;
mem[16'h9A70] = 8'h42;
mem[16'h9A71] = 8'h46;
mem[16'h9A72] = 8'h4A;
mem[16'h9A73] = 8'h52;
mem[16'h9A74] = 8'h62;
mem[16'h9A75] = 8'h42;
mem[16'h9A76] = 8'h42;
mem[16'h9A77] = 8'h00;
mem[16'h9A78] = 8'h3C;
mem[16'h9A79] = 8'h42;
mem[16'h9A7A] = 8'h42;
mem[16'h9A7B] = 8'h42;
mem[16'h9A7C] = 8'h42;
mem[16'h9A7D] = 8'h42;
mem[16'h9A7E] = 8'h3C;
mem[16'h9A7F] = 8'h00;
mem[16'h9A80] = 8'h3E;
mem[16'h9A81] = 8'h42;
mem[16'h9A82] = 8'h42;
mem[16'h9A83] = 8'h3E;
mem[16'h9A84] = 8'h02;
mem[16'h9A85] = 8'h02;
mem[16'h9A86] = 8'h02;
mem[16'h9A87] = 8'h00;
mem[16'h9A88] = 8'h3C;
mem[16'h9A89] = 8'h42;
mem[16'h9A8A] = 8'h42;
mem[16'h9A8B] = 8'h42;
mem[16'h9A8C] = 8'h52;
mem[16'h9A8D] = 8'h22;
mem[16'h9A8E] = 8'h5C;
mem[16'h9A8F] = 8'h00;
mem[16'h9A90] = 8'h3E;
mem[16'h9A91] = 8'h42;
mem[16'h9A92] = 8'h42;
mem[16'h9A93] = 8'h3E;
mem[16'h9A94] = 8'h12;
mem[16'h9A95] = 8'h22;
mem[16'h9A96] = 8'h42;
mem[16'h9A97] = 8'h00;
mem[16'h9A98] = 8'h3C;
mem[16'h9A99] = 8'h42;
mem[16'h9A9A] = 8'h02;
mem[16'h9A9B] = 8'h3C;
mem[16'h9A9C] = 8'h40;
mem[16'h9A9D] = 8'h42;
mem[16'h9A9E] = 8'h3C;
mem[16'h9A9F] = 8'h00;
mem[16'h9AA0] = 8'h7C;
mem[16'h9AA1] = 8'h10;
mem[16'h9AA2] = 8'h10;
mem[16'h9AA3] = 8'h10;
mem[16'h9AA4] = 8'h10;
mem[16'h9AA5] = 8'h10;
mem[16'h9AA6] = 8'h10;
mem[16'h9AA7] = 8'h00;
mem[16'h9AA8] = 8'h42;
mem[16'h9AA9] = 8'h42;
mem[16'h9AAA] = 8'h42;
mem[16'h9AAB] = 8'h42;
mem[16'h9AAC] = 8'h42;
mem[16'h9AAD] = 8'h42;
mem[16'h9AAE] = 8'h3C;
mem[16'h9AAF] = 8'h00;
mem[16'h9AB0] = 8'h42;
mem[16'h9AB1] = 8'h42;
mem[16'h9AB2] = 8'h42;
mem[16'h9AB3] = 8'h24;
mem[16'h9AB4] = 8'h24;
mem[16'h9AB5] = 8'h18;
mem[16'h9AB6] = 8'h18;
mem[16'h9AB7] = 8'h00;
mem[16'h9AB8] = 8'h42;
mem[16'h9AB9] = 8'h42;
mem[16'h9ABA] = 8'h42;
mem[16'h9ABB] = 8'h5A;
mem[16'h9ABC] = 8'h5A;
mem[16'h9ABD] = 8'h66;
mem[16'h9ABE] = 8'h42;
mem[16'h9ABF] = 8'h00;
mem[16'h9AC0] = 8'h42;
mem[16'h9AC1] = 8'h42;
mem[16'h9AC2] = 8'h24;
mem[16'h9AC3] = 8'h18;
mem[16'h9AC4] = 8'h24;
mem[16'h9AC5] = 8'h42;
mem[16'h9AC6] = 8'h42;
mem[16'h9AC7] = 8'h00;
mem[16'h9AC8] = 8'h44;
mem[16'h9AC9] = 8'h44;
mem[16'h9ACA] = 8'h44;
mem[16'h9ACB] = 8'h38;
mem[16'h9ACC] = 8'h10;
mem[16'h9ACD] = 8'h10;
mem[16'h9ACE] = 8'h10;
mem[16'h9ACF] = 8'h00;
mem[16'h9AD0] = 8'h7E;
mem[16'h9AD1] = 8'h40;
mem[16'h9AD2] = 8'h20;
mem[16'h9AD3] = 8'h18;
mem[16'h9AD4] = 8'h04;
mem[16'h9AD5] = 8'h02;
mem[16'h9AD6] = 8'h7E;
mem[16'h9AD7] = 8'h00;
mem[16'h9AD8] = 8'h3C;
mem[16'h9AD9] = 8'h04;
mem[16'h9ADA] = 8'h04;
mem[16'h9ADB] = 8'h04;
mem[16'h9ADC] = 8'h04;
mem[16'h9ADD] = 8'h04;
mem[16'h9ADE] = 8'h3C;
mem[16'h9ADF] = 8'h00;
mem[16'h9AE0] = 8'h00;
mem[16'h9AE1] = 8'h02;
mem[16'h9AE2] = 8'h04;
mem[16'h9AE3] = 8'h08;
mem[16'h9AE4] = 8'h10;
mem[16'h9AE5] = 8'h20;
mem[16'h9AE6] = 8'h40;
mem[16'h9AE7] = 8'h00;
mem[16'h9AE8] = 8'h3C;
mem[16'h9AE9] = 8'h20;
mem[16'h9AEA] = 8'h20;
mem[16'h9AEB] = 8'h20;
mem[16'h9AEC] = 8'h20;
mem[16'h9AED] = 8'h20;
mem[16'h9AEE] = 8'h3C;
mem[16'h9AEF] = 8'h00;
mem[16'h9AF0] = 8'h10;
mem[16'h9AF1] = 8'h28;
mem[16'h9AF2] = 8'h44;
mem[16'h9AF3] = 8'h00;
mem[16'h9AF4] = 8'h00;
mem[16'h9AF5] = 8'h00;
mem[16'h9AF6] = 8'h00;
mem[16'h9AF7] = 8'h00;
mem[16'h9AF8] = 8'h02;
mem[16'h9AF9] = 8'h00;
mem[16'h9AFA] = 8'h00;
mem[16'h9AFB] = 8'h00;
mem[16'h9AFC] = 8'h00;
mem[16'h9AFD] = 8'h00;
mem[16'h9AFE] = 8'h00;
mem[16'h9AFF] = 8'hFF;
mem[16'h9B00] = 8'h08;
mem[16'h9B01] = 8'h10;
mem[16'h9B02] = 8'h20;
mem[16'h9B03] = 8'h00;
mem[16'h9B04] = 8'h00;
mem[16'h9B05] = 8'h00;
mem[16'h9B06] = 8'h00;
mem[16'h9B07] = 8'h00;
mem[16'h9B08] = 8'h00;
mem[16'h9B09] = 8'h00;
mem[16'h9B0A] = 8'h1C;
mem[16'h9B0B] = 8'h20;
mem[16'h9B0C] = 8'h3C;
mem[16'h9B0D] = 8'h22;
mem[16'h9B0E] = 8'h5C;
mem[16'h9B0F] = 8'h00;
mem[16'h9B10] = 8'h02;
mem[16'h9B11] = 8'h02;
mem[16'h9B12] = 8'h3A;
mem[16'h9B13] = 8'h46;
mem[16'h9B14] = 8'h42;
mem[16'h9B15] = 8'h46;
mem[16'h9B16] = 8'h3A;
mem[16'h9B17] = 8'h00;
mem[16'h9B18] = 8'h00;
mem[16'h9B19] = 8'h00;
mem[16'h9B1A] = 8'h3C;
mem[16'h9B1B] = 8'h02;
mem[16'h9B1C] = 8'h02;
mem[16'h9B1D] = 8'h02;
mem[16'h9B1E] = 8'h3C;
mem[16'h9B1F] = 8'h00;
mem[16'h9B20] = 8'h40;
mem[16'h9B21] = 8'h40;
mem[16'h9B22] = 8'h5C;
mem[16'h9B23] = 8'h62;
mem[16'h9B24] = 8'h42;
mem[16'h9B25] = 8'h62;
mem[16'h9B26] = 8'h5C;
mem[16'h9B27] = 8'h00;
mem[16'h9B28] = 8'h00;
mem[16'h9B29] = 8'h00;
mem[16'h9B2A] = 8'h3C;
mem[16'h9B2B] = 8'h42;
mem[16'h9B2C] = 8'h7E;
mem[16'h9B2D] = 8'h02;
mem[16'h9B2E] = 8'h3C;
mem[16'h9B2F] = 8'h00;
mem[16'h9B30] = 8'h30;
mem[16'h9B31] = 8'h48;
mem[16'h9B32] = 8'h08;
mem[16'h9B33] = 8'h3E;
mem[16'h9B34] = 8'h08;
mem[16'h9B35] = 8'h08;
mem[16'h9B36] = 8'h08;
mem[16'h9B37] = 8'h00;
mem[16'h9B38] = 8'h00;
mem[16'h9B39] = 8'h00;
mem[16'h9B3A] = 8'h5C;
mem[16'h9B3B] = 8'h62;
mem[16'h9B3C] = 8'h62;
mem[16'h9B3D] = 8'h5C;
mem[16'h9B3E] = 8'h40;
mem[16'h9B3F] = 8'h3C;
mem[16'h9B40] = 8'h02;
mem[16'h9B41] = 8'h02;
mem[16'h9B42] = 8'h3A;
mem[16'h9B43] = 8'h46;
mem[16'h9B44] = 8'h42;
mem[16'h9B45] = 8'h42;
mem[16'h9B46] = 8'h42;
mem[16'h9B47] = 8'h00;
mem[16'h9B48] = 8'h10;
mem[16'h9B49] = 8'h00;
mem[16'h9B4A] = 8'h18;
mem[16'h9B4B] = 8'h10;
mem[16'h9B4C] = 8'h10;
mem[16'h9B4D] = 8'h10;
mem[16'h9B4E] = 8'h38;
mem[16'h9B4F] = 8'h00;
mem[16'h9B50] = 8'h20;
mem[16'h9B51] = 8'h00;
mem[16'h9B52] = 8'h30;
mem[16'h9B53] = 8'h20;
mem[16'h9B54] = 8'h20;
mem[16'h9B55] = 8'h20;
mem[16'h9B56] = 8'h22;
mem[16'h9B57] = 8'h1C;
mem[16'h9B58] = 8'h02;
mem[16'h9B59] = 8'h02;
mem[16'h9B5A] = 8'h22;
mem[16'h9B5B] = 8'h12;
mem[16'h9B5C] = 8'h0A;
mem[16'h9B5D] = 8'h16;
mem[16'h9B5E] = 8'h22;
mem[16'h9B5F] = 8'h00;
mem[16'h9B60] = 8'h18;
mem[16'h9B61] = 8'h10;
mem[16'h9B62] = 8'h10;
mem[16'h9B63] = 8'h10;
mem[16'h9B64] = 8'h10;
mem[16'h9B65] = 8'h10;
mem[16'h9B66] = 8'h38;
mem[16'h9B67] = 8'h00;
mem[16'h9B68] = 8'h00;
mem[16'h9B69] = 8'h00;
mem[16'h9B6A] = 8'h2E;
mem[16'h9B6B] = 8'h54;
mem[16'h9B6C] = 8'h54;
mem[16'h9B6D] = 8'h54;
mem[16'h9B6E] = 8'h54;
mem[16'h9B6F] = 8'h00;
mem[16'h9B70] = 8'h00;
mem[16'h9B71] = 8'h00;
mem[16'h9B72] = 8'h3E;
mem[16'h9B73] = 8'h44;
mem[16'h9B74] = 8'h44;
mem[16'h9B75] = 8'h44;
mem[16'h9B76] = 8'h44;
mem[16'h9B77] = 8'h00;
mem[16'h9B78] = 8'h00;
mem[16'h9B79] = 8'h00;
mem[16'h9B7A] = 8'h38;
mem[16'h9B7B] = 8'h44;
mem[16'h9B7C] = 8'h44;
mem[16'h9B7D] = 8'h44;
mem[16'h9B7E] = 8'h38;
mem[16'h9B7F] = 8'h00;
mem[16'h9B80] = 8'h00;
mem[16'h9B81] = 8'h00;
mem[16'h9B82] = 8'h3A;
mem[16'h9B83] = 8'h46;
mem[16'h9B84] = 8'h46;
mem[16'h9B85] = 8'h3A;
mem[16'h9B86] = 8'h02;
mem[16'h9B87] = 8'h02;
mem[16'h9B88] = 8'h00;
mem[16'h9B89] = 8'h00;
mem[16'h9B8A] = 8'h5C;
mem[16'h9B8B] = 8'h62;
mem[16'h9B8C] = 8'h62;
mem[16'h9B8D] = 8'h5C;
mem[16'h9B8E] = 8'h40;
mem[16'h9B8F] = 8'h40;
mem[16'h9B90] = 8'h00;
mem[16'h9B91] = 8'h00;
mem[16'h9B92] = 8'h3A;
mem[16'h9B93] = 8'h46;
mem[16'h9B94] = 8'h02;
mem[16'h9B95] = 8'h02;
mem[16'h9B96] = 8'h02;
mem[16'h9B97] = 8'h00;
mem[16'h9B98] = 8'h00;
mem[16'h9B99] = 8'h00;
mem[16'h9B9A] = 8'h7C;
mem[16'h9B9B] = 8'h02;
mem[16'h9B9C] = 8'h3C;
mem[16'h9B9D] = 8'h40;
mem[16'h9B9E] = 8'h3E;
mem[16'h9B9F] = 8'h00;
mem[16'h9BA0] = 8'h08;
mem[16'h9BA1] = 8'h08;
mem[16'h9BA2] = 8'h3E;
mem[16'h9BA3] = 8'h08;
mem[16'h9BA4] = 8'h08;
mem[16'h9BA5] = 8'h48;
mem[16'h9BA6] = 8'h30;
mem[16'h9BA7] = 8'h00;
mem[16'h9BA8] = 8'h00;
mem[16'h9BA9] = 8'h00;
mem[16'h9BAA] = 8'h42;
mem[16'h9BAB] = 8'h42;
mem[16'h9BAC] = 8'h42;
mem[16'h9BAD] = 8'h62;
mem[16'h9BAE] = 8'h5C;
mem[16'h9BAF] = 8'h00;
mem[16'h9BB0] = 8'h00;
mem[16'h9BB1] = 8'h00;
mem[16'h9BB2] = 8'h42;
mem[16'h9BB3] = 8'h42;
mem[16'h9BB4] = 8'h42;
mem[16'h9BB5] = 8'h24;
mem[16'h9BB6] = 8'h18;
mem[16'h9BB7] = 8'h00;
mem[16'h9BB8] = 8'h00;
mem[16'h9BB9] = 8'h00;
mem[16'h9BBA] = 8'h44;
mem[16'h9BBB] = 8'h44;
mem[16'h9BBC] = 8'h54;
mem[16'h9BBD] = 8'h54;
mem[16'h9BBE] = 8'h6C;
mem[16'h9BBF] = 8'h00;
mem[16'h9BC0] = 8'h00;
mem[16'h9BC1] = 8'h00;
mem[16'h9BC2] = 8'h42;
mem[16'h9BC3] = 8'h24;
mem[16'h9BC4] = 8'h18;
mem[16'h9BC5] = 8'h24;
mem[16'h9BC6] = 8'h42;
mem[16'h9BC7] = 8'h00;
mem[16'h9BC8] = 8'h00;
mem[16'h9BC9] = 8'h00;
mem[16'h9BCA] = 8'h42;
mem[16'h9BCB] = 8'h42;
mem[16'h9BCC] = 8'h62;
mem[16'h9BCD] = 8'h5C;
mem[16'h9BCE] = 8'h40;
mem[16'h9BCF] = 8'h3C;
mem[16'h9BD0] = 8'h00;
mem[16'h9BD1] = 8'h00;
mem[16'h9BD2] = 8'h7E;
mem[16'h9BD3] = 8'h20;
mem[16'h9BD4] = 8'h18;
mem[16'h9BD5] = 8'h04;
mem[16'h9BD6] = 8'h7E;
mem[16'h9BD7] = 8'h00;
mem[16'h9BD8] = 8'h38;
mem[16'h9BD9] = 8'h04;
mem[16'h9BDA] = 8'h04;
mem[16'h9BDB] = 8'h06;
mem[16'h9BDC] = 8'h04;
mem[16'h9BDD] = 8'h04;
mem[16'h9BDE] = 8'h38;
mem[16'h9BDF] = 8'h00;
mem[16'h9BE0] = 8'h08;
mem[16'h9BE1] = 8'h08;
mem[16'h9BE2] = 8'h08;
mem[16'h9BE3] = 8'h08;
mem[16'h9BE4] = 8'h08;
mem[16'h9BE5] = 8'h08;
mem[16'h9BE6] = 8'h08;
mem[16'h9BE7] = 8'h08;
mem[16'h9BE8] = 8'h0E;
mem[16'h9BE9] = 8'h10;
mem[16'h9BEA] = 8'h10;
mem[16'h9BEB] = 8'h30;
mem[16'h9BEC] = 8'h10;
mem[16'h9BED] = 8'h10;
mem[16'h9BEE] = 8'h0E;
mem[16'h9BEF] = 8'h00;
mem[16'h9BF0] = 8'h28;
mem[16'h9BF1] = 8'h14;
mem[16'h9BF2] = 8'h00;
mem[16'h9BF3] = 8'h00;
mem[16'h9BF4] = 8'h00;
mem[16'h9BF5] = 8'h00;
mem[16'h9BF6] = 8'h00;
mem[16'h9BF7] = 8'h00;
mem[16'h9BF8] = 8'hFF;
mem[16'h9BF9] = 8'hFF;
mem[16'h9BFA] = 8'hFF;
mem[16'h9BFB] = 8'hFF;
mem[16'h9BFC] = 8'hFF;
mem[16'h9BFD] = 8'h0F;
mem[16'h9BFE] = 8'hAB;
mem[16'h9BFF] = 8'h81;
mem[16'h9C00] = 8'h4C;
mem[16'h9C01] = 8'h5F;
mem[16'h9C02] = 8'h9C;
mem[16'h9C03] = 8'hA9;
mem[16'h9C04] = 8'h00;
mem[16'h9C05] = 8'h8D;
mem[16'h9C06] = 8'h06;
mem[16'h9C07] = 8'hA0;
mem[16'h9C08] = 8'h8D;
mem[16'h9C09] = 8'h09;
mem[16'h9C0A] = 8'hA0;
mem[16'h9C0B] = 8'h8D;
mem[16'h9C0C] = 8'h0A;
mem[16'h9C0D] = 8'hA0;
mem[16'h9C0E] = 8'hA9;
mem[16'h9C0F] = 8'h05;
mem[16'h9C10] = 8'h8D;
mem[16'h9C11] = 8'h07;
mem[16'h9C12] = 8'hA0;
mem[16'h9C13] = 8'hAD;
mem[16'h9C14] = 8'h19;
mem[16'h9C15] = 8'hA0;
mem[16'h9C16] = 8'hC9;
mem[16'h9C17] = 8'h1F;
mem[16'h9C18] = 8'hD0;
mem[16'h9C19] = 8'h1A;
mem[16'h9C1A] = 8'h10;
mem[16'h9C1B] = 8'h01;
mem[16'h9C1C] = 8'h85;
mem[16'h9C1D] = 8'hCD;
mem[16'h9C1E] = 8'h10;
mem[16'h9C1F] = 8'hC0;
mem[16'h9C20] = 8'hCE;
mem[16'h9C21] = 8'hF3;
mem[16'h9C22] = 8'h03;
mem[16'h9C23] = 8'hD0;
mem[16'h9C24] = 8'hFB;
mem[16'h9C25] = 8'hAD;
mem[16'h9C26] = 8'h00;
mem[16'h9C27] = 8'hC0;
mem[16'h9C28] = 8'h30;
mem[16'h9C29] = 8'h0A;
mem[16'h9C2A] = 8'hCE;
mem[16'h9C2B] = 8'hF4;
mem[16'h9C2C] = 8'h03;
mem[16'h9C2D] = 8'hD0;
mem[16'h9C2E] = 8'hF1;
mem[16'h9C2F] = 8'hCE;
mem[16'h9C30] = 8'h19;
mem[16'h9C31] = 8'hA0;
mem[16'h9C32] = 8'hD0;
mem[16'h9C33] = 8'hEC;
mem[16'h9C34] = 8'hA9;
mem[16'h9C35] = 8'h1F;
mem[16'h9C36] = 8'h8D;
mem[16'h9C37] = 8'h19;
mem[16'h9C38] = 8'hA0;
mem[16'h9C39] = 8'h20;
mem[16'h9C3A] = 8'h00;
mem[16'h9C3B] = 8'h0D;
mem[16'h9C3C] = 8'hEA;
mem[16'h9C3D] = 8'hEA;
mem[16'h9C3E] = 8'hA9;
mem[16'h9C3F] = 8'hFF;
mem[16'h9C40] = 8'h85;
mem[16'h9C41] = 8'h3A;
mem[16'h9C42] = 8'hA9;
mem[16'h9C43] = 8'hBF;
mem[16'h9C44] = 8'h85;
mem[16'h9C45] = 8'h3B;
mem[16'h9C46] = 8'hA0;
mem[16'h9C47] = 8'h13;
mem[16'h9C48] = 8'hD1;
mem[16'h9C49] = 8'h3A;
mem[16'h9C4A] = 8'hA0;
mem[16'h9C4B] = 8'h07;
mem[16'h9C4C] = 8'hB1;
mem[16'h9C4D] = 8'h3A;
mem[16'h9C4E] = 8'hC9;
mem[16'h9C4F] = 8'hA0;
mem[16'h9C50] = 8'hD0;
mem[16'h9C51] = 8'h02;
mem[16'h9C52] = 8'h60;
mem[16'h9C53] = 8'hA9;
mem[16'h9C54] = 8'hC9;
mem[16'h9C55] = 8'hC4;
mem[16'h9C56] = 8'hF0;
mem[16'h9C57] = 8'hFA;
mem[16'h9C58] = 8'hC9;
mem[16'h9C59] = 8'hCA;
mem[16'h9C5A] = 8'hF0;
mem[16'h9C5B] = 8'hF6;
mem[16'h9C5C] = 8'h4C;
mem[16'h9C5D] = 8'h4A;
mem[16'h9C5E] = 8'h9C;
mem[16'h9C5F] = 8'hA0;
mem[16'h9C60] = 8'h00;
mem[16'h9C61] = 8'h84;
mem[16'h9C62] = 8'h00;
mem[16'h9C63] = 8'h84;
mem[16'h9C64] = 8'h02;
mem[16'h9C65] = 8'hA9;
mem[16'h9C66] = 8'h97;
mem[16'h9C67] = 8'h85;
mem[16'h9C68] = 8'h01;
mem[16'h9C69] = 8'hA9;
mem[16'h9C6A] = 8'h03;
mem[16'h9C6B] = 8'h85;
mem[16'h9C6C] = 8'h03;
mem[16'h9C6D] = 8'hA2;
mem[16'h9C6E] = 8'h05;
mem[16'h9C6F] = 8'hAD;
mem[16'h9C70] = 8'h55;
mem[16'h9C71] = 8'hC0;
mem[16'h9C72] = 8'hEA;
mem[16'h9C73] = 8'hEA;
mem[16'h9C74] = 8'hEA;
mem[16'h9C75] = 8'hEA;
mem[16'h9C76] = 8'hEA;
mem[16'h9C77] = 8'hEA;
mem[16'h9C78] = 8'hEA;
mem[16'h9C79] = 8'hEA;
mem[16'h9C7A] = 8'hEA;
mem[16'h9C7B] = 8'hB1;
mem[16'h9C7C] = 8'h00;
mem[16'h9C7D] = 8'h91;
mem[16'h9C7E] = 8'h02;
mem[16'h9C7F] = 8'hC8;
mem[16'h9C80] = 8'hD0;
mem[16'h9C81] = 8'hF9;
mem[16'h9C82] = 8'hE6;
mem[16'h9C83] = 8'h01;
mem[16'h9C84] = 8'hE6;
mem[16'h9C85] = 8'h03;
mem[16'h9C86] = 8'hCA;
mem[16'h9C87] = 8'hD0;
mem[16'h9C88] = 8'hF2;
mem[16'h9C89] = 8'h4C;
mem[16'h9C8A] = 8'h03;
mem[16'h9C8B] = 8'h40;
mem[16'h9C8C] = 8'h84;
mem[16'h9C8D] = 8'hC2;
mem[16'h9C8E] = 8'hCC;
mem[16'h9C8F] = 8'hCF;
mem[16'h9C90] = 8'hED;
mem[16'h9C91] = 8'hFD;
mem[16'h9C92] = 8'h20;
mem[16'h9C93] = 8'h3A;
mem[16'h9C94] = 8'hFF;
mem[16'h9C95] = 8'hA9;
mem[16'h9C96] = 8'hA1;
mem[16'h9C97] = 8'h85;
mem[16'h9C98] = 8'h33;
mem[16'h9C99] = 8'h20;
mem[16'h9C9A] = 8'h67;
mem[16'h9C9B] = 8'hFD;
mem[16'h9C9C] = 8'h20;
mem[16'h9C9D] = 8'hC7;
mem[16'h9C9E] = 8'hFF;
mem[16'h9C9F] = 8'hAD;
mem[16'h9CA0] = 8'h00;
mem[16'h9CA1] = 8'h02;
mem[16'h9CA2] = 8'hC9;
mem[16'h9CA3] = 8'hA0;
mem[16'h9CA4] = 8'hF0;
mem[16'h9CA5] = 8'h13;
mem[16'h9CA6] = 8'hC8;
mem[16'h9CA7] = 8'hC9;
mem[16'h9CA8] = 8'hA4;
mem[16'h9CA9] = 8'hF0;
mem[16'h9CAA] = 8'h92;
mem[16'h9CAB] = 8'h88;
mem[16'h9CAC] = 8'h20;
mem[16'h9CAD] = 8'hA7;
mem[16'h9CAE] = 8'hFF;
mem[16'h9CAF] = 8'hC9;
mem[16'h9CB0] = 8'h93;
mem[16'h9CB1] = 8'hD0;
mem[16'h9CB2] = 8'hD5;
mem[16'h9CB3] = 8'h8A;
mem[16'h9CB4] = 8'hF0;
mem[16'h9CB5] = 8'hD2;
mem[16'h9CB6] = 8'h20;
mem[16'h9CB7] = 8'h78;
mem[16'h9CB8] = 8'hFE;
mem[16'h9CB9] = 8'hA9;
mem[16'h9CBA] = 8'h03;
mem[16'h9CBB] = 8'h85;
mem[16'h9CBC] = 8'h3D;
mem[16'h9CBD] = 8'h20;
mem[16'h9CBE] = 8'h34;
mem[16'h9CBF] = 8'hF6;
mem[16'h9CC0] = 8'h0A;
mem[16'h9CC1] = 8'hE9;
mem[16'h9CC2] = 8'hBE;
mem[16'h9CC3] = 8'hC9;
mem[16'h9CC4] = 8'hC2;
mem[16'h9CC5] = 8'h90;
mem[16'h9CC6] = 8'hC1;
mem[16'h9CC7] = 8'h0A;
mem[16'h9CC8] = 8'h0A;
mem[16'h9CC9] = 8'hA2;
mem[16'h9CCA] = 8'h04;
mem[16'h9CCB] = 8'h0A;
mem[16'h9CCC] = 8'h26;
mem[16'h9CCD] = 8'h42;
mem[16'h9CCE] = 8'h26;
mem[16'h9CCF] = 8'h43;
mem[16'h9CD0] = 8'hCA;
mem[16'h9CD1] = 8'h10;
mem[16'h9CD2] = 8'hF8;
mem[16'h9CD3] = 8'hC6;
mem[16'h9CD4] = 8'h3D;
mem[16'h9CD5] = 8'hF0;
mem[16'h9CD6] = 8'hF4;
mem[16'h9CD7] = 8'h10;
mem[16'h9CD8] = 8'hE4;
mem[16'h9CD9] = 8'hA2;
mem[16'h9CDA] = 8'h05;
mem[16'h9CDB] = 8'h20;
mem[16'h9CDC] = 8'h34;
mem[16'h9CDD] = 8'hF6;
mem[16'h9CDE] = 8'h84;
mem[16'h9CDF] = 8'h34;
mem[16'h9CE0] = 8'hDD;
mem[16'h9CE1] = 8'hB4;
mem[16'h9CE2] = 8'hF9;
mem[16'h9CE3] = 8'hD0;
mem[16'h9CE4] = 8'h13;
mem[16'h9CE5] = 8'h20;
mem[16'h9CE6] = 8'h34;
mem[16'h9CE7] = 8'hF6;
mem[16'h9CE8] = 8'hDD;
mem[16'h9CE9] = 8'hBA;
mem[16'h9CEA] = 8'hF9;
mem[16'h9CEB] = 8'hF0;
mem[16'h9CEC] = 8'h0D;
mem[16'h9CED] = 8'hBD;
mem[16'h9CEE] = 8'hBA;
mem[16'h9CEF] = 8'hF9;
mem[16'h9CF0] = 8'hF0;
mem[16'h9CF1] = 8'h07;
mem[16'h9CF2] = 8'hC9;
mem[16'h9CF3] = 8'hA4;
mem[16'h9CF4] = 8'hF0;
mem[16'h9CF5] = 8'h03;
mem[16'h9CF6] = 8'hA4;
mem[16'h9CF7] = 8'h34;
mem[16'h9CF8] = 8'h18;
mem[16'h9CF9] = 8'h88;
mem[16'h9CFA] = 8'h26;
mem[16'h9CFB] = 8'h44;
mem[16'h9CFC] = 8'hE0;
mem[16'h9CFD] = 8'h03;
mem[16'h9CFE] = 8'hD0;
mem[16'h9CFF] = 8'h0D;
mem[16'h9D00] = 8'hB3;
mem[16'h9D01] = 8'hBD;
mem[16'h9D02] = 8'hC8;
mem[16'h9D03] = 8'hB4;
mem[16'h9D04] = 8'h29;
mem[16'h9D05] = 8'h7F;
mem[16'h9D06] = 8'h0D;
mem[16'h9D07] = 8'h9E;
mem[16'h9D08] = 8'hB3;
mem[16'h9D09] = 8'h9D;
mem[16'h9D0A] = 8'hC8;
mem[16'h9D0B] = 8'hB4;
mem[16'h9D0C] = 8'h20;
mem[16'h9D0D] = 8'h37;
mem[16'h9D0E] = 8'hB0;
mem[16'h9D0F] = 8'h4C;
mem[16'h9D10] = 8'h7F;
mem[16'h9D11] = 8'hB3;
mem[16'h9D12] = 8'h20;
mem[16'h9D13] = 8'h00;
mem[16'h9D14] = 8'hB3;
mem[16'h9D15] = 8'h4C;
mem[16'h9D16] = 8'h7F;
mem[16'h9D17] = 8'hB3;
mem[16'h9D18] = 8'h20;
mem[16'h9D19] = 8'h28;
mem[16'h9D1A] = 8'hAB;
mem[16'h9D1B] = 8'h20;
mem[16'h9D1C] = 8'hB6;
mem[16'h9D1D] = 8'hB0;
mem[16'h9D1E] = 8'hB0;
mem[16'h9D1F] = 8'hEF;
mem[16'h9D20] = 8'hEE;
mem[16'h9D21] = 8'hE4;
mem[16'h9D22] = 8'hB5;
mem[16'h9D23] = 8'hD0;
mem[16'h9D24] = 8'hF6;
mem[16'h9D25] = 8'hEE;
mem[16'h9D26] = 8'hE5;
mem[16'h9D27] = 8'hB5;
mem[16'h9D28] = 8'h4C;
mem[16'h9D29] = 8'h1B;
mem[16'h9D2A] = 8'hAD;
mem[16'h9D2B] = 8'h20;
mem[16'h9D2C] = 8'h28;
mem[16'h9D2D] = 8'hAB;
mem[16'h9D2E] = 8'hAE;
mem[16'h9D2F] = 8'h9C;
mem[16'h9D30] = 8'hB3;
mem[16'h9D31] = 8'hBD;
mem[16'h9D32] = 8'hC8;
mem[16'h9D33] = 8'hB4;
mem[16'h9D34] = 8'h10;
mem[16'h9D35] = 8'h03;
mem[16'h9D36] = 8'h4C;
mem[16'h9D37] = 8'h7B;
mem[16'h9D38] = 8'hB3;
mem[16'h9D39] = 8'hAE;
mem[16'h9D3A] = 8'h9C;
mem[16'h9D3B] = 8'hB3;
mem[16'h9D3C] = 8'hBD;
mem[16'h9D3D] = 8'hC6;
mem[16'h9D3E] = 8'hB4;
mem[16'h9D3F] = 8'h8D;
mem[16'h9D40] = 8'hD1;
mem[16'h9D41] = 8'hB5;
mem[16'h9D42] = 8'h9D;
mem[16'h9D43] = 8'hE6;
mem[16'h9D44] = 8'hB4;
mem[16'h9D45] = 8'hA9;
mem[16'h9D46] = 8'hFF;
mem[16'h9D47] = 8'h9D;
mem[16'h9D48] = 8'hC6;
mem[16'h9D49] = 8'hB4;
mem[16'h9D4A] = 8'hBC;
mem[16'h9D4B] = 8'hC7;
mem[16'h9D4C] = 8'hB4;
mem[16'h9D4D] = 8'h8C;
mem[16'h9D4E] = 8'hD2;
mem[16'h9D4F] = 8'hB5;
mem[16'h9D50] = 8'h20;
mem[16'h9D51] = 8'h37;
mem[16'h9D52] = 8'hB0;
mem[16'h9D53] = 8'h18;
mem[16'h9D54] = 8'h20;
mem[16'h9D55] = 8'h5E;
mem[16'h9D56] = 8'hAF;
mem[16'h9D57] = 8'hB0;
mem[16'h9D58] = 8'h2A;
mem[16'h9D59] = 8'h20;
mem[16'h9D5A] = 8'h0C;
mem[16'h9D5B] = 8'hAF;
mem[16'h9D5C] = 8'hA0;
mem[16'h9D5D] = 8'h0C;
mem[16'h9D5E] = 8'h8C;
mem[16'h9D5F] = 8'h9C;
mem[16'h9D60] = 8'hB3;
mem[16'h9D61] = 8'hB1;
mem[16'h9D62] = 8'h42;
mem[16'h9D63] = 8'h30;
mem[16'h9D64] = 8'h0B;
mem[16'h9D65] = 8'hF0;
mem[16'h9D66] = 8'h09;
mem[16'h9D67] = 8'h48;
mem[16'h9D68] = 8'hC8;
mem[16'h9D69] = 8'hB1;
mem[16'h9D6A] = 8'h42;
mem[16'h9D6B] = 8'hA8;
mem[16'h9D6C] = 8'h68;
mem[16'h9D6D] = 8'h20;
mem[16'h9D6E] = 8'h89;
mem[16'h9D6F] = 8'hAD;
mem[16'h9D70] = 8'hAC;
mem[16'h9D71] = 8'h9C;
mem[16'h9D72] = 8'hB3;
mem[16'h9D73] = 8'hC8;
mem[16'h9D74] = 8'hC8;
mem[16'h9D75] = 8'hD0;
mem[16'h9D76] = 8'hE7;
mem[16'h9D77] = 8'hAD;
mem[16'h9D78] = 8'hD3;
mem[16'h9D79] = 8'hB5;
mem[16'h9D7A] = 8'hAC;
mem[16'h9D7B] = 8'hD4;
mem[16'h9D7C] = 8'hB5;
mem[16'h9D7D] = 8'h20;
mem[16'h9D7E] = 8'h89;
mem[16'h9D7F] = 8'hAD;
mem[16'h9D80] = 8'h38;
mem[16'h9D81] = 8'hB0;
mem[16'h9D82] = 8'hD1;
mem[16'h9D83] = 8'h20;
mem[16'h9D84] = 8'hFB;
mem[16'h9D85] = 8'hAF;
mem[16'h9D86] = 8'h4C;
mem[16'h9D87] = 8'h7F;
mem[16'h9D88] = 8'hB3;
mem[16'h9D89] = 8'h38;
mem[16'h9D8A] = 8'h20;
mem[16'h9D8B] = 8'hDD;
mem[16'h9D8C] = 8'hB2;
mem[16'h9D8D] = 8'hA9;
mem[16'h9D8E] = 8'h00;
mem[16'h9D8F] = 8'hA2;
mem[16'h9D90] = 8'h05;
mem[16'h9D91] = 8'h9D;
mem[16'h9D92] = 8'hF0;
mem[16'h9D93] = 8'hB5;
mem[16'h9D94] = 8'hCA;
mem[16'h9D95] = 8'h10;
mem[16'h9D96] = 8'hFA;
mem[16'h9D97] = 8'h60;
mem[16'h9D98] = 8'h20;
mem[16'h9D99] = 8'hDC;
mem[16'h9D9A] = 8'hAB;
mem[16'h9D9B] = 8'hA9;
mem[16'h9D9C] = 8'hFF;
mem[16'h9D9D] = 8'h8D;
mem[16'h9D9E] = 8'hF9;
mem[16'h9D9F] = 8'hB5;
mem[16'h9DA0] = 8'h20;
mem[16'h9DA1] = 8'hF7;
mem[16'h9DA2] = 8'hAF;
mem[16'h9DA3] = 8'hA9;
mem[16'h9DA4] = 8'h16;
mem[16'h9DA5] = 8'h8D;
mem[16'h9DA6] = 8'h9D;
mem[16'h9DA7] = 8'hB3;
mem[16'h9DA8] = 8'h20;
mem[16'h9DA9] = 8'h2F;
mem[16'h9DAA] = 8'hAE;
mem[16'h9DAB] = 8'h20;
mem[16'h9DAC] = 8'h2F;
mem[16'h9DAD] = 8'hAE;
mem[16'h9DAE] = 8'hA2;
mem[16'h9DAF] = 8'h0B;
mem[16'h9DB0] = 8'hBD;
mem[16'h9DB1] = 8'hAF;
mem[16'h9DB2] = 8'hB3;
mem[16'h9DB3] = 8'h20;
mem[16'h9DB4] = 8'hED;
mem[16'h9DB5] = 8'hFD;
mem[16'h9DB6] = 8'hCA;
mem[16'h9DB7] = 8'h10;
mem[16'h9DB8] = 8'hF7;
mem[16'h9DB9] = 8'h86;
mem[16'h9DBA] = 8'h45;
mem[16'h9DBB] = 8'hAD;
mem[16'h9DBC] = 8'hF6;
mem[16'h9DBD] = 8'hB7;
mem[16'h9DBE] = 8'h85;
mem[16'h9DBF] = 8'h44;
mem[16'h9DC0] = 8'h20;
mem[16'h9DC1] = 8'h42;
mem[16'h9DC2] = 8'hAE;
mem[16'h9DC3] = 8'h20;
mem[16'h9DC4] = 8'h2F;
mem[16'h9DC5] = 8'hAE;
mem[16'h9DC6] = 8'h20;
mem[16'h9DC7] = 8'h2F;
mem[16'h9DC8] = 8'hAE;
mem[16'h9DC9] = 8'h18;
mem[16'h9DCA] = 8'h20;
mem[16'h9DCB] = 8'h11;
mem[16'h9DCC] = 8'hB0;
mem[16'h9DCD] = 8'hB0;
mem[16'h9DCE] = 8'h5D;
mem[16'h9DCF] = 8'hA2;
mem[16'h9DD0] = 8'h00;
mem[16'h9DD1] = 8'h8E;
mem[16'h9DD2] = 8'h9C;
mem[16'h9DD3] = 8'hB3;
mem[16'h9DD4] = 8'hBD;
mem[16'h9DD5] = 8'hC6;
mem[16'h9DD6] = 8'hB4;
mem[16'h9DD7] = 8'hF0;
mem[16'h9DD8] = 8'h53;
mem[16'h9DD9] = 8'h30;
mem[16'h9DDA] = 8'h4A;
mem[16'h9DDB] = 8'hA0;
mem[16'h9DDC] = 8'hA0;
mem[16'h9DDD] = 8'hBD;
mem[16'h9DDE] = 8'hC8;
mem[16'h9DDF] = 8'hB4;
mem[16'h9DE0] = 8'h10;
mem[16'h9DE1] = 8'h02;
mem[16'h9DE2] = 8'hA0;
mem[16'h9DE3] = 8'hAA;
mem[16'h9DE4] = 8'h98;
mem[16'h9DE5] = 8'h20;
mem[16'h9DE6] = 8'hED;
mem[16'h9DE7] = 8'hFD;
mem[16'h9DE8] = 8'hBD;
mem[16'h9DE9] = 8'hC8;
mem[16'h9DEA] = 8'hB4;
mem[16'h9DEB] = 8'h29;
mem[16'h9DEC] = 8'h7F;
mem[16'h9DED] = 8'hA0;
mem[16'h9DEE] = 8'h07;
mem[16'h9DEF] = 8'h0A;
mem[16'h9DF0] = 8'h0A;
mem[16'h9DF1] = 8'hB0;
mem[16'h9DF2] = 8'h03;
mem[16'h9DF3] = 8'h88;
mem[16'h9DF4] = 8'hD0;
mem[16'h9DF5] = 8'hFA;
mem[16'h9DF6] = 8'hB9;
mem[16'h9DF7] = 8'hA7;
mem[16'h9DF8] = 8'hB3;
mem[16'h9DF9] = 8'h20;
mem[16'h9DFA] = 8'hED;
mem[16'h9DFB] = 8'hFD;
mem[16'h9DFC] = 8'hA9;
mem[16'h9DFD] = 8'hA0;
mem[16'h9DFE] = 8'h20;
mem[16'h9DFF] = 8'hED;
mem[16'h9E00] = 8'hFD;
mem[16'h9E01] = 8'hBD;
mem[16'h9E02] = 8'hE7;
mem[16'h9E03] = 8'hB4;
mem[16'h9E04] = 8'h85;
mem[16'h9E05] = 8'h44;
mem[16'h9E06] = 8'hBD;
mem[16'h9E07] = 8'hE8;
mem[16'h9E08] = 8'hB4;
mem[16'h9E09] = 8'h85;
mem[16'h9E0A] = 8'h45;
mem[16'h9E0B] = 8'h20;
mem[16'h9E0C] = 8'h42;
mem[16'h9E0D] = 8'hAE;
mem[16'h9E0E] = 8'hA9;
mem[16'h9E0F] = 8'hA0;
mem[16'h9E10] = 8'h20;
mem[16'h9E11] = 8'hED;
mem[16'h9E12] = 8'hFD;
mem[16'h9E13] = 8'hE8;
mem[16'h9E14] = 8'hE8;
mem[16'h9E15] = 8'hE8;
mem[16'h9E16] = 8'hA0;
mem[16'h9E17] = 8'h1D;
mem[16'h9E18] = 8'hBD;
mem[16'h9E19] = 8'hC6;
mem[16'h9E1A] = 8'hB4;
mem[16'h9E1B] = 8'h20;
mem[16'h9E1C] = 8'hED;
mem[16'h9E1D] = 8'hFD;
mem[16'h9E1E] = 8'hE8;
mem[16'h9E1F] = 8'h88;
mem[16'h9E20] = 8'h10;
mem[16'h9E21] = 8'hF6;
mem[16'h9E22] = 8'h20;
mem[16'h9E23] = 8'h2F;
mem[16'h9E24] = 8'hAE;
mem[16'h9E25] = 8'h20;
mem[16'h9E26] = 8'h30;
mem[16'h9E27] = 8'hB2;
mem[16'h9E28] = 8'h90;
mem[16'h9E29] = 8'hA7;
mem[16'h9E2A] = 8'hB0;
mem[16'h9E2B] = 8'h9E;
mem[16'h9E2C] = 8'h4C;
mem[16'h9E2D] = 8'h7F;
mem[16'h9E2E] = 8'hB3;
mem[16'h9E2F] = 8'hA9;
mem[16'h9E30] = 8'h8D;
mem[16'h9E31] = 8'h20;
mem[16'h9E32] = 8'hED;
mem[16'h9E33] = 8'hFD;
mem[16'h9E34] = 8'hCE;
mem[16'h9E35] = 8'h9D;
mem[16'h9E36] = 8'hB3;
mem[16'h9E37] = 8'hD0;
mem[16'h9E38] = 8'h08;
mem[16'h9E39] = 8'h20;
mem[16'h9E3A] = 8'h0C;
mem[16'h9E3B] = 8'hFD;
mem[16'h9E3C] = 8'hA9;
mem[16'h9E3D] = 8'h15;
mem[16'h9E3E] = 8'h8D;
mem[16'h9E3F] = 8'h9D;
mem[16'h9E40] = 8'hB3;
mem[16'h9E41] = 8'h60;
mem[16'h9E42] = 8'hA0;
mem[16'h9E43] = 8'h02;
mem[16'h9E44] = 8'hA9;
mem[16'h9E45] = 8'h00;
mem[16'h9E46] = 8'h48;
mem[16'h9E47] = 8'hA5;
mem[16'h9E48] = 8'h44;
mem[16'h9E49] = 8'hD9;
mem[16'h9E4A] = 8'hA4;
mem[16'h9E4B] = 8'hB3;
mem[16'h9E4C] = 8'h90;
mem[16'h9E4D] = 8'h12;
mem[16'h9E4E] = 8'hF9;
mem[16'h9E4F] = 8'hA4;
mem[16'h9E50] = 8'hB3;
mem[16'h9E51] = 8'h85;
mem[16'h9E52] = 8'h44;
mem[16'h9E53] = 8'hA5;
mem[16'h9E54] = 8'h45;
mem[16'h9E55] = 8'hE9;
mem[16'h9E56] = 8'h00;
mem[16'h9E57] = 8'h85;
mem[16'h9E58] = 8'h45;
mem[16'h9E59] = 8'h68;
mem[16'h9E5A] = 8'h69;
mem[16'h9E5B] = 8'h00;
mem[16'h9E5C] = 8'h48;
mem[16'h9E5D] = 8'h4C;
mem[16'h9E5E] = 8'h47;
mem[16'h9E5F] = 8'hAE;
mem[16'h9E60] = 8'h68;
mem[16'h9E61] = 8'h09;
mem[16'h9E62] = 8'hB0;
mem[16'h9E63] = 8'h20;
mem[16'h9E64] = 8'hED;
mem[16'h9E65] = 8'hFD;
mem[16'h9E66] = 8'h88;
mem[16'h9E67] = 8'h10;
mem[16'h9E68] = 8'hDB;
mem[16'h9E69] = 8'h60;
mem[16'h9E6A] = 8'h20;
mem[16'h9E6B] = 8'h08;
mem[16'h9E6C] = 8'hAF;
mem[16'h9E6D] = 8'hA0;
mem[16'h9E6E] = 8'h00;
mem[16'h9E6F] = 8'h8C;
mem[16'h9E70] = 8'hC5;
mem[16'h9E71] = 8'hB5;
mem[16'h9E72] = 8'hB1;
mem[16'h9E73] = 8'h42;
mem[16'h9E74] = 8'h99;
mem[16'h9E75] = 8'hD1;
mem[16'h9E76] = 8'hB5;
mem[16'h9E77] = 8'hC8;
mem[16'h9E78] = 8'hC0;
mem[16'h9E79] = 8'h2D;
mem[16'h9E7A] = 8'hD0;
mem[16'h9E7B] = 8'hF6;
mem[16'h9E7C] = 8'h18;
mem[16'h9E7D] = 8'h60;
mem[16'h9E7E] = 8'h20;
mem[16'h9E7F] = 8'h08;
mem[16'h9E80] = 8'hAF;
mem[16'h9E81] = 8'hA0;
mem[16'h9E82] = 8'h00;
mem[16'h9E83] = 8'hB9;
mem[16'h9E84] = 8'hD1;
mem[16'h9E85] = 8'hB5;
mem[16'h9E86] = 8'h91;
mem[16'h9E87] = 8'h42;
mem[16'h9E88] = 8'hC8;
mem[16'h9E89] = 8'hC0;
mem[16'h9E8A] = 8'h2D;
mem[16'h9E8B] = 8'hD0;
mem[16'h9E8C] = 8'hF6;
mem[16'h9E8D] = 8'h60;
mem[16'h9E8E] = 8'h20;
mem[16'h9E8F] = 8'hDC;
mem[16'h9E90] = 8'hAB;
mem[16'h9E91] = 8'hA9;
mem[16'h9E92] = 8'h04;
mem[16'h9E93] = 8'h20;
mem[16'h9E94] = 8'h58;
mem[16'h9E95] = 8'hB0;
mem[16'h9E96] = 8'hAD;
mem[16'h9E97] = 8'hF9;
mem[16'h9E98] = 8'hB5;
mem[16'h9E99] = 8'h49;
mem[16'h9E9A] = 8'hFF;
mem[16'h9E9B] = 8'h8D;
mem[16'h9E9C] = 8'hC1;
mem[16'h9E9D] = 8'hB3;
mem[16'h9E9E] = 8'hA9;
mem[16'h9E9F] = 8'h11;
mem[16'h9EA0] = 8'h8D;
mem[16'h9EA1] = 8'hEB;
mem[16'h9EA2] = 8'hB3;
mem[16'h9EA3] = 8'hA9;
mem[16'h9EA4] = 8'h01;
mem[16'h9EA5] = 8'h8D;
mem[16'h9EA6] = 8'hEC;
mem[16'h9EA7] = 8'hB3;
mem[16'h9EA8] = 8'hA2;
mem[16'h9EA9] = 8'h38;
mem[16'h9EAA] = 8'hA9;
mem[16'h9EAB] = 8'h00;
mem[16'h9EAC] = 8'h9D;
mem[16'h9EAD] = 8'hBB;
mem[16'h9EAE] = 8'hB3;
mem[16'h9EAF] = 8'hE8;
mem[16'h9EB0] = 8'hD0;
mem[16'h9EB1] = 8'hFA;
mem[16'h9EB2] = 8'hA2;
mem[16'h9EB3] = 8'h0C;
mem[16'h9EB4] = 8'hE0;
mem[16'h9EB5] = 8'h8C;
mem[16'h9EB6] = 8'hF0;
mem[16'h9EB7] = 8'h14;
mem[16'h9EB8] = 8'hA0;
mem[16'h9EB9] = 8'h03;
mem[16'h9EBA] = 8'hB9;
mem[16'h9EBB] = 8'hA0;
mem[16'h9EBC] = 8'hB3;
mem[16'h9EBD] = 8'h9D;
mem[16'h9EBE] = 8'hF3;
mem[16'h9EBF] = 8'hB3;
mem[16'h9EC0] = 8'hE8;
mem[16'h9EC1] = 8'h88;
mem[16'h9EC2] = 8'h10;
mem[16'h9EC3] = 8'hF6;
mem[16'h9EC4] = 8'hE0;
mem[16'h9EC5] = 8'h44;
mem[16'h9EC6] = 8'hD0;
mem[16'h9EC7] = 8'hEC;
mem[16'h9EC8] = 8'hA2;
mem[16'h9EC9] = 8'h48;
mem[16'h9ECA] = 8'hD0;
mem[16'h9ECB] = 8'hE8;
mem[16'h9ECC] = 8'h20;
mem[16'h9ECD] = 8'hFB;
mem[16'h9ECE] = 8'hAF;
mem[16'h9ECF] = 8'hA2;
mem[16'h9ED0] = 8'h00;
mem[16'h9ED1] = 8'h8A;
mem[16'h9ED2] = 8'h9D;
mem[16'h9ED3] = 8'hBB;
mem[16'h9ED4] = 8'hB4;
mem[16'h9ED5] = 8'hE8;
mem[16'h9ED6] = 8'hD0;
mem[16'h9ED7] = 8'hFA;
mem[16'h9ED8] = 8'h20;
mem[16'h9ED9] = 8'h45;
mem[16'h9EDA] = 8'hB0;
mem[16'h9EDB] = 8'hA9;
mem[16'h9EDC] = 8'h11;
mem[16'h9EDD] = 8'hAC;
mem[16'h9EDE] = 8'hF0;
mem[16'h9EDF] = 8'hB3;
mem[16'h9EE0] = 8'h88;
mem[16'h9EE1] = 8'h88;
mem[16'h9EE2] = 8'h8D;
mem[16'h9EE3] = 8'hEC;
mem[16'h9EE4] = 8'hB7;
mem[16'h9EE5] = 8'h8D;
mem[16'h9EE6] = 8'hBC;
mem[16'h9EE7] = 8'hB4;
mem[16'h9EE8] = 8'h8C;
mem[16'h9EE9] = 8'hBD;
mem[16'h9EEA] = 8'hB4;
mem[16'h9EEB] = 8'hC8;
mem[16'h9EEC] = 8'h8C;
mem[16'h9EED] = 8'hED;
mem[16'h9EEE] = 8'hB7;
mem[16'h9EEF] = 8'hA9;
mem[16'h9EF0] = 8'h02;
mem[16'h9EF1] = 8'h20;
mem[16'h9EF2] = 8'h58;
mem[16'h9EF3] = 8'hB0;
mem[16'h9EF4] = 8'hAC;
mem[16'h9EF5] = 8'hBD;
mem[16'h9EF6] = 8'hB4;
mem[16'h9EF7] = 8'h88;
mem[16'h9EF8] = 8'h30;
mem[16'h9EF9] = 8'h05;
mem[16'h9EFA] = 8'hD0;
mem[16'h9EFB] = 8'hEC;
mem[16'h9EFC] = 8'h98;
mem[16'h9EFD] = 8'hF0;
mem[16'h9EFE] = 8'hE6;
mem[16'h9EFF] = 8'h20;
mem[16'h9F00] = 8'hC2;
mem[16'h9F01] = 8'hB7;
mem[16'h9F02] = 8'h20;
mem[16'h9F03] = 8'h4A;
mem[16'h9F04] = 8'hB7;
mem[16'h9F05] = 8'h4C;
mem[16'h9F06] = 8'h7F;
mem[16'h9F07] = 8'hB3;
mem[16'h9F08] = 8'hA2;
mem[16'h9F09] = 8'h00;
mem[16'h9F0A] = 8'hF0;
mem[16'h9F0B] = 8'h06;
mem[16'h9F0C] = 8'hA2;
mem[16'h9F0D] = 8'h02;
mem[16'h9F0E] = 8'hD0;
mem[16'h9F0F] = 8'h02;
mem[16'h9F10] = 8'hA2;
mem[16'h9F11] = 8'h04;
mem[16'h9F12] = 8'hBD;
mem[16'h9F13] = 8'hC7;
mem[16'h9F14] = 8'hB5;
mem[16'h9F15] = 8'h85;
mem[16'h9F16] = 8'h42;
mem[16'h9F17] = 8'hBD;
mem[16'h9F18] = 8'hC8;
mem[16'h9F19] = 8'hB5;
mem[16'h9F1A] = 8'h85;
mem[16'h9F1B] = 8'h43;
mem[16'h9F1C] = 8'h60;
mem[16'h9F1D] = 8'h2C;
mem[16'h9F1E] = 8'hD5;
mem[16'h9F1F] = 8'hB5;
mem[16'h9F20] = 8'h70;
mem[16'h9F21] = 8'h01;
mem[16'h9F22] = 8'h60;
mem[16'h9F23] = 8'h20;
mem[16'h9F24] = 8'hE4;
mem[16'h9F25] = 8'hAF;
mem[16'h9F26] = 8'hA9;
mem[16'h9F27] = 8'h02;
mem[16'h9F28] = 8'h20;
mem[16'h9F29] = 8'h52;
mem[16'h9F2A] = 8'hB0;
mem[16'h9F2B] = 8'hA9;
mem[16'h9F2C] = 8'hBF;
mem[16'h9F2D] = 8'h2D;
mem[16'h9F2E] = 8'hD5;
mem[16'h9F2F] = 8'hB5;
mem[16'h9F30] = 8'h8D;
mem[16'h9F31] = 8'hD5;
mem[16'h9F32] = 8'hB5;
mem[16'h9F33] = 8'h60;
mem[16'h9F34] = 8'hAD;
mem[16'h9F35] = 8'hD5;
mem[16'h9F36] = 8'hB5;
mem[16'h9F37] = 8'h30;
mem[16'h9F38] = 8'h01;
mem[16'h9F39] = 8'h60;
mem[16'h9F3A] = 8'h20;
mem[16'h9F3B] = 8'h4B;
mem[16'h9F3C] = 8'hAF;
mem[16'h9F3D] = 8'hA9;
mem[16'h9F3E] = 8'h02;
mem[16'h9F3F] = 8'h20;
mem[16'h9F40] = 8'h52;
mem[16'h9F41] = 8'hB0;
mem[16'h9F42] = 8'hA9;
mem[16'h9F43] = 8'h7F;
mem[16'h9F44] = 8'h2D;
mem[16'h9F45] = 8'hD5;
mem[16'h9F46] = 8'hB5;
mem[16'h9F47] = 8'h8D;
mem[16'h9F48] = 8'hD5;
mem[16'h9F49] = 8'hB5;
mem[16'h9F4A] = 8'h60;
mem[16'h9F4B] = 8'hAD;
mem[16'h9F4C] = 8'hC9;
mem[16'h9F4D] = 8'hB5;
mem[16'h9F4E] = 8'h8D;
mem[16'h9F4F] = 8'hF0;
mem[16'h9F50] = 8'hB7;
mem[16'h9F51] = 8'hAD;
mem[16'h9F52] = 8'hCA;
mem[16'h9F53] = 8'hB5;
mem[16'h9F54] = 8'h8D;
mem[16'h9F55] = 8'hF1;
mem[16'h9F56] = 8'hB7;
mem[16'h9F57] = 8'hAE;
mem[16'h9F58] = 8'hD3;
mem[16'h9F59] = 8'hB5;
mem[16'h9F5A] = 8'hAC;
mem[16'h9F5B] = 8'hD4;
mem[16'h9F5C] = 8'hB5;
mem[16'h9F5D] = 8'h60;
mem[16'h9F5E] = 8'h08;
mem[16'h9F5F] = 8'h20;
mem[16'h9F60] = 8'h34;
mem[16'h9F61] = 8'hAF;
mem[16'h9F62] = 8'h20;
mem[16'h9F63] = 8'h4B;
mem[16'h9F64] = 8'hAF;
mem[16'h9F65] = 8'h20;
mem[16'h9F66] = 8'h0C;
mem[16'h9F67] = 8'hAF;
mem[16'h9F68] = 8'h28;
mem[16'h9F69] = 8'hB0;
mem[16'h9F6A] = 8'h09;
mem[16'h9F6B] = 8'hAE;
mem[16'h9F6C] = 8'hD1;
mem[16'h9F6D] = 8'hB5;
mem[16'h9F6E] = 8'hAC;
mem[16'h9F6F] = 8'hD2;
mem[16'h9F70] = 8'hB5;
mem[16'h9F71] = 8'h4C;
mem[16'h9F72] = 8'hB5;
mem[16'h9F73] = 8'hAF;
mem[16'h9F74] = 8'hA0;
mem[16'h9F75] = 8'h01;
mem[16'h9F76] = 8'hB1;
mem[16'h9F77] = 8'h42;
mem[16'h9F78] = 8'hF0;
mem[16'h9F79] = 8'h08;
mem[16'h9F7A] = 8'hAA;
mem[16'h9F7B] = 8'hC8;
mem[16'h9F7C] = 8'hB1;
mem[16'h9F7D] = 8'h42;
mem[16'h9F7E] = 8'hA8;
mem[16'h9F7F] = 8'h4C;
mem[16'h9F80] = 8'hB5;
mem[16'h9F81] = 8'hAF;
mem[16'h9F82] = 8'hAD;
mem[16'h9F83] = 8'hBB;
mem[16'h9F84] = 8'hB5;
mem[16'h9F85] = 8'hC9;
mem[16'h9F86] = 8'h04;
mem[16'h9F87] = 8'hF0;
mem[16'h9F88] = 8'h02;
mem[16'h9F89] = 8'h38;
mem[16'h9F8A] = 8'h60;
mem[16'h9F8B] = 8'h20;
mem[16'h9F8C] = 8'h44;
mem[16'h9F8D] = 8'hB2;
mem[16'h9F8E] = 8'hA0;
mem[16'h9F8F] = 8'h02;
mem[16'h9F90] = 8'h91;
mem[16'h9F91] = 8'h42;
mem[16'h9F92] = 8'h48;
mem[16'h9F93] = 8'h88;
mem[16'h9F94] = 8'hAD;
mem[16'h9F95] = 8'hF1;
mem[16'h9F96] = 8'hB5;
mem[16'h9F97] = 8'h91;
mem[16'h9F98] = 8'h42;
mem[16'h9F99] = 8'h48;
mem[16'h9F9A] = 8'h20;
mem[16'h9F9B] = 8'h3A;
mem[16'h9F9C] = 8'hAF;
mem[16'h9F9D] = 8'h20;
mem[16'h9F9E] = 8'hD6;
mem[16'h9F9F] = 8'hB7;
mem[16'h9FA0] = 8'hA0;
mem[16'h9FA1] = 8'h05;
mem[16'h9FA2] = 8'hAD;
mem[16'h9FA3] = 8'hDE;
mem[16'h9FA4] = 8'hB5;
mem[16'h9FA5] = 8'h91;
mem[16'h9FA6] = 8'h42;
mem[16'h9FA7] = 8'hC8;
mem[16'h9FA8] = 8'hAD;
mem[16'h9FA9] = 8'hDF;
mem[16'h9FAA] = 8'hB5;
mem[16'h9FAB] = 8'h91;
mem[16'h9FAC] = 8'h42;
mem[16'h9FAD] = 8'h68;
mem[16'h9FAE] = 8'hAA;
mem[16'h9FAF] = 8'h68;
mem[16'h9FB0] = 8'hA8;
mem[16'h9FB1] = 8'hA9;
mem[16'h9FB2] = 8'h02;
mem[16'h9FB3] = 8'hD0;
mem[16'h9FB4] = 8'h02;
mem[16'h9FB5] = 8'hA9;
mem[16'h9FB6] = 8'h01;
mem[16'h9FB7] = 8'h8E;
mem[16'h9FB8] = 8'hD3;
mem[16'h9FB9] = 8'hB5;
mem[16'h9FBA] = 8'h8C;
mem[16'h9FBB] = 8'hD4;
mem[16'h9FBC] = 8'hB5;
mem[16'h9FBD] = 8'h20;
mem[16'h9FBE] = 8'h52;
mem[16'h9FBF] = 8'hB0;
mem[16'h9FC0] = 8'hA0;
mem[16'h9FC1] = 8'h05;
mem[16'h9FC2] = 8'hB1;
mem[16'h9FC3] = 8'h42;
mem[16'h9FC4] = 8'h8D;
mem[16'h9FC5] = 8'hDC;
mem[16'h9FC6] = 8'hB5;
mem[16'h9FC7] = 8'h18;
mem[16'h9FC8] = 8'h6D;
mem[16'h9FC9] = 8'hDA;
mem[16'h9FCA] = 8'hB5;
mem[16'h9FCB] = 8'h8D;
mem[16'h9FCC] = 8'hDE;
mem[16'h9FCD] = 8'hB5;
mem[16'h9FCE] = 8'hC8;
mem[16'h9FCF] = 8'hB1;
mem[16'h9FD0] = 8'h42;
mem[16'h9FD1] = 8'h8D;
mem[16'h9FD2] = 8'hDD;
mem[16'h9FD3] = 8'hB5;
mem[16'h9FD4] = 8'h6D;
mem[16'h9FD5] = 8'hDB;
mem[16'h9FD6] = 8'hB5;
mem[16'h9FD7] = 8'h8D;
mem[16'h9FD8] = 8'hDF;
mem[16'h9FD9] = 8'hB5;
mem[16'h9FDA] = 8'h18;
mem[16'h9FDB] = 8'h60;
mem[16'h9FDC] = 8'h20;
mem[16'h9FDD] = 8'hE4;
mem[16'h9FDE] = 8'hAF;
mem[16'h9FDF] = 8'hA9;
mem[16'h9FE0] = 8'h01;
mem[16'h9FE1] = 8'h4C;
mem[16'h9FE2] = 8'h52;
mem[16'h9FE3] = 8'hB0;
mem[16'h9FE4] = 8'hAC;
mem[16'h9FE5] = 8'hCB;
mem[16'h9FE6] = 8'hB5;
mem[16'h9FE7] = 8'hAD;
mem[16'h9FE8] = 8'hCC;
mem[16'h9FE9] = 8'hB5;
mem[16'h9FEA] = 8'h8C;
mem[16'h9FEB] = 8'hF0;
mem[16'h9FEC] = 8'hB7;
mem[16'h9FED] = 8'h8D;
mem[16'h9FEE] = 8'hF1;
mem[16'h9FEF] = 8'hB7;
mem[16'h9FF0] = 8'hAE;
mem[16'h9FF1] = 8'hD6;
mem[16'h9FF2] = 8'hB5;
mem[16'h9FF3] = 8'hAC;
mem[16'h9FF4] = 8'hD7;
mem[16'h9FF5] = 8'hB5;
mem[16'h9FF6] = 8'h60;
mem[16'h9FF7] = 8'hA9;
mem[16'h9FF8] = 8'h01;
mem[16'h9FF9] = 8'hD0;
mem[16'h9FFA] = 8'h02;
mem[16'h9FFB] = 8'hA9;
mem[16'h9FFC] = 8'h02;
mem[16'h9FFD] = 8'hAC;
mem[16'h9FFE] = 8'hC3;
mem[16'h9FFF] = 8'hAA;
mem[16'hA000] = 8'h0B;
mem[16'hA001] = 8'h60;
mem[16'hA002] = 8'h01;
mem[16'hA003] = 8'hCD;
mem[16'hA004] = 8'hB2;
mem[16'hA005] = 8'hAA;
mem[16'hA006] = 8'h00;
mem[16'hA007] = 8'h05;
mem[16'hA008] = 8'h00;
mem[16'hA009] = 8'h00;
mem[16'hA00A] = 8'h00;
mem[16'hA00B] = 8'hAD;
mem[16'hA00C] = 8'h01;
mem[16'hA00D] = 8'h02;
mem[16'hA00E] = 8'hC9;
mem[16'hA00F] = 8'h8D;
mem[16'hA010] = 8'h41;
mem[16'hA011] = 8'h00;
mem[16'hA012] = 8'h00;
mem[16'hA013] = 8'h00;
mem[16'hA014] = 8'h00;
mem[16'hA015] = 8'h00;
mem[16'hA016] = 8'hBE;
mem[16'hA017] = 8'h00;
mem[16'hA018] = 8'h4C;
mem[16'hA019] = 8'h1F;
mem[16'hA01A] = 8'h60;
mem[16'hA01B] = 8'h00;
mem[16'hA01C] = 8'hFF;
mem[16'hA01D] = 8'hAA;
mem[16'hA01E] = 8'hAC;
mem[16'hA01F] = 8'h5F;
mem[16'hA020] = 8'hAA;
mem[16'hA021] = 8'h20;
mem[16'hA022] = 8'h5E;
mem[16'hA023] = 8'hA6;
mem[16'hA024] = 8'h90;
mem[16'hA025] = 8'h0C;
mem[16'hA026] = 8'hA9;
mem[16'hA027] = 8'h02;
mem[16'hA028] = 8'h39;
mem[16'hA029] = 8'h09;
mem[16'hA02A] = 8'hA9;
mem[16'hA02B] = 8'hF0;
mem[16'hA02C] = 8'h05;
mem[16'hA02D] = 8'hA9;
mem[16'hA02E] = 8'h0F;
mem[16'hA02F] = 8'h4C;
mem[16'hA030] = 8'hD2;
mem[16'hA031] = 8'hA6;
mem[16'hA032] = 8'hC0;
mem[16'hA033] = 8'h06;
mem[16'hA034] = 8'hD0;
mem[16'hA035] = 8'h02;
mem[16'hA036] = 8'h84;
mem[16'hA037] = 8'h33;
mem[16'hA038] = 8'hA9;
mem[16'hA039] = 8'h20;
mem[16'hA03A] = 8'h39;
mem[16'hA03B] = 8'h09;
mem[16'hA03C] = 8'hA9;
mem[16'hA03D] = 8'hF0;
mem[16'hA03E] = 8'h61;
mem[16'hA03F] = 8'h20;
mem[16'hA040] = 8'h95;
mem[16'hA041] = 8'hA0;
mem[16'hA042] = 8'h08;
mem[16'hA043] = 8'h20;
mem[16'hA044] = 8'hA4;
mem[16'hA045] = 8'hA1;
mem[16'hA046] = 8'hF0;
mem[16'hA047] = 8'h1E;
mem[16'hA048] = 8'h0A;
mem[16'hA049] = 8'h90;
mem[16'hA04A] = 8'h05;
mem[16'hA04B] = 8'h30;
mem[16'hA04C] = 8'h03;
mem[16'hA04D] = 8'h4C;
mem[16'hA04E] = 8'h00;
mem[16'hA04F] = 8'hA0;
mem[16'hA050] = 8'h6A;
mem[16'hA051] = 8'h4C;
mem[16'hA052] = 8'h59;
mem[16'hA053] = 8'hA0;
mem[16'hA054] = 8'h20;
mem[16'hA055] = 8'h93;
mem[16'hA056] = 8'hA1;
mem[16'hA057] = 8'hF0;
mem[16'hA058] = 8'h0D;
mem[16'hA059] = 8'h99;
mem[16'hA05A] = 8'h75;
mem[16'hA05B] = 8'hAA;
mem[16'hA05C] = 8'hC8;
mem[16'hA05D] = 8'hC0;
mem[16'hA05E] = 8'h3C;
mem[16'hA05F] = 8'h90;
mem[16'hA060] = 8'hF3;
mem[16'hA061] = 8'h20;
mem[16'hA062] = 8'h93;
mem[16'hA063] = 8'hA1;
mem[16'hA064] = 8'hD0;
mem[16'hA065] = 8'hFB;
mem[16'hA066] = 8'h28;
mem[16'hA067] = 8'hD0;
mem[16'hA068] = 8'h0F;
mem[16'hA069] = 8'hAC;
mem[16'hA06A] = 8'h5F;
mem[16'hA06B] = 8'hAA;
mem[16'hA06C] = 8'hA9;
mem[16'hA06D] = 8'h10;
mem[16'hA06E] = 8'h39;
mem[16'hA06F] = 8'h09;
mem[16'hA070] = 8'hA9;
mem[16'hA071] = 8'hF0;
mem[16'hA072] = 8'h0C;
mem[16'hA073] = 8'hA0;
mem[16'hA074] = 8'h1E;
mem[16'hA075] = 8'h08;
mem[16'hA076] = 8'hD0;
mem[16'hA077] = 8'hCB;
mem[16'hA078] = 8'hAD;
mem[16'hA079] = 8'h93;
mem[16'hA07A] = 8'hAA;
mem[16'hA07B] = 8'hC9;
mem[16'hA07C] = 8'hA0;
mem[16'hA07D] = 8'hF0;
mem[16'hA07E] = 8'h13;
mem[16'hA07F] = 8'hAD;
mem[16'hA080] = 8'h75;
mem[16'hA081] = 8'hAA;
mem[16'hA082] = 8'hC9;
mem[16'hA083] = 8'hA0;
mem[16'hA084] = 8'hD0;
mem[16'hA085] = 8'h4B;
mem[16'hA086] = 8'hAC;
mem[16'hA087] = 8'h5F;
mem[16'hA088] = 8'hAA;
mem[16'hA089] = 8'hA9;
mem[16'hA08A] = 8'hC0;
mem[16'hA08B] = 8'h39;
mem[16'hA08C] = 8'h09;
mem[16'hA08D] = 8'hA9;
mem[16'hA08E] = 8'hF0;
mem[16'hA08F] = 8'h02;
mem[16'hA090] = 8'h10;
mem[16'hA091] = 8'h3F;
mem[16'hA092] = 8'h4C;
mem[16'hA093] = 8'h00;
mem[16'hA094] = 8'hA0;
mem[16'hA095] = 8'hA0;
mem[16'hA096] = 8'h3C;
mem[16'hA097] = 8'hA9;
mem[16'hA098] = 8'hA0;
mem[16'hA099] = 8'h99;
mem[16'hA09A] = 8'h74;
mem[16'hA09B] = 8'hAA;
mem[16'hA09C] = 8'h88;
mem[16'hA09D] = 8'hD0;
mem[16'hA09E] = 8'hFA;
mem[16'hA09F] = 8'h60;
mem[16'hA0A0] = 8'h8D;
mem[16'hA0A1] = 8'h75;
mem[16'hA0A2] = 8'hAA;
mem[16'hA0A3] = 8'hA9;
mem[16'hA0A4] = 8'h0C;
mem[16'hA0A5] = 8'h39;
mem[16'hA0A6] = 8'h09;
mem[16'hA0A7] = 8'hA9;
mem[16'hA0A8] = 8'hF0;
mem[16'hA0A9] = 8'h27;
mem[16'hA0AA] = 8'h20;
mem[16'hA0AB] = 8'hB9;
mem[16'hA0AC] = 8'hA1;
mem[16'hA0AD] = 8'hB0;
mem[16'hA0AE] = 8'h1F;
mem[16'hA0AF] = 8'hA8;
mem[16'hA0B0] = 8'hD0;
mem[16'hA0B1] = 8'h17;
mem[16'hA0B2] = 8'hE0;
mem[16'hA0B3] = 8'h11;
mem[16'hA0B4] = 8'hB0;
mem[16'hA0B5] = 8'h13;
mem[16'hA0B6] = 8'hAC;
mem[16'hA0B7] = 8'h5F;
mem[16'hA0B8] = 8'hAA;
mem[16'hA0B9] = 8'hA9;
mem[16'hA0BA] = 8'h08;
mem[16'hA0BB] = 8'h39;
mem[16'hA0BC] = 8'h09;
mem[16'hA0BD] = 8'hA9;
mem[16'hA0BE] = 8'hF0;
mem[16'hA0BF] = 8'h06;
mem[16'hA0C0] = 8'hE0;
mem[16'hA0C1] = 8'h08;
mem[16'hA0C2] = 8'hB0;
mem[16'hA0C3] = 8'hCE;
mem[16'hA0C4] = 8'h90;
mem[16'hA0C5] = 8'h0B;
mem[16'hA0C6] = 8'h8A;
mem[16'hA0C7] = 8'hD0;
mem[16'hA0C8] = 8'h08;
mem[16'hA0C9] = 8'hA9;
mem[16'hA0CA] = 8'h02;
mem[16'hA0CB] = 8'h4C;
mem[16'hA0CC] = 8'hD2;
mem[16'hA0CD] = 8'hA6;
mem[16'hA0CE] = 8'h4C;
mem[16'hA0CF] = 8'hC4;
mem[16'hA0D0] = 8'hA6;
mem[16'hA0D1] = 8'hA9;
mem[16'hA0D2] = 8'h00;
mem[16'hA0D3] = 8'h8D;
mem[16'hA0D4] = 8'h65;
mem[16'hA0D5] = 8'hAA;
mem[16'hA0D6] = 8'h8D;
mem[16'hA0D7] = 8'h74;
mem[16'hA0D8] = 8'hAA;
mem[16'hA0D9] = 8'h8D;
mem[16'hA0DA] = 8'h66;
mem[16'hA0DB] = 8'hAA;
mem[16'hA0DC] = 8'h8D;
mem[16'hA0DD] = 8'h6C;
mem[16'hA0DE] = 8'hAA;
mem[16'hA0DF] = 8'h8D;
mem[16'hA0E0] = 8'h6D;
mem[16'hA0E1] = 8'hAA;
mem[16'hA0E2] = 8'h20;
mem[16'hA0E3] = 8'hDC;
mem[16'hA0E4] = 8'hBF;
mem[16'hA0E5] = 8'hAD;
mem[16'hA0E6] = 8'h5D;
mem[16'hA0E7] = 8'hAA;
mem[16'hA0E8] = 8'h20;
mem[16'hA0E9] = 8'hA4;
mem[16'hA0EA] = 8'hA1;
mem[16'hA0EB] = 8'hD0;
mem[16'hA0EC] = 8'h1F;
mem[16'hA0ED] = 8'hC9;
mem[16'hA0EE] = 8'h8D;
mem[16'hA0EF] = 8'hD0;
mem[16'hA0F0] = 8'hF7;
mem[16'hA0F1] = 8'hAE;
mem[16'hA0F2] = 8'h5F;
mem[16'hA0F3] = 8'hAA;
mem[16'hA0F4] = 8'hAD;
mem[16'hA0F5] = 8'h65;
mem[16'hA0F6] = 8'hAA;
mem[16'hA0F7] = 8'h1D;
mem[16'hA0F8] = 8'h0A;
mem[16'hA0F9] = 8'hA9;
mem[16'hA0FA] = 8'h5D;
mem[16'hA0FB] = 8'h0A;
mem[16'hA0FC] = 8'hA9;
mem[16'hA0FD] = 8'hD0;
mem[16'hA0FE] = 8'h93;
mem[16'hA0FF] = 8'hAE;
mem[16'hA100] = 8'h00;
mem[16'hA101] = 8'hAA;
mem[16'hA102] = 8'h00;
mem[16'hA103] = 8'h76;
mem[16'hA104] = 8'h00;
mem[16'hA105] = 8'h63;
mem[16'hA106] = 8'h00;
mem[16'hA107] = 8'h8E;
mem[16'hA108] = 8'h00;
mem[16'hA109] = 8'hAA;
mem[16'hA10A] = 8'h00;
mem[16'hA10B] = 8'hDC;
mem[16'hA10C] = 8'h00;
mem[16'hA10D] = 8'h0A;
mem[16'hA10E] = 8'h00;
mem[16'hA10F] = 8'h40;
mem[16'hA110] = 8'h00;
mem[16'hA111] = 8'hF0;
mem[16'hA112] = 8'h00;
mem[16'hA113] = 8'hCA;
mem[16'hA114] = 8'h00;
mem[16'hA115] = 8'hF8;
mem[16'hA116] = 8'h00;
mem[16'hA117] = 8'hB6;
mem[16'hA118] = 8'h00;
mem[16'hA119] = 8'h4A;
mem[16'hA11A] = 8'h00;
mem[16'hA11B] = 8'h30;
mem[16'hA11C] = 8'h00;
mem[16'hA11D] = 8'h0D;
mem[16'hA11E] = 8'h00;
mem[16'hA11F] = 8'hAA;
mem[16'hA120] = 8'h00;
mem[16'hA121] = 8'h65;
mem[16'hA122] = 8'h00;
mem[16'hA123] = 8'hCA;
mem[16'hA124] = 8'h00;
mem[16'hA125] = 8'h64;
mem[16'hA126] = 8'h00;
mem[16'hA127] = 8'h20;
mem[16'hA128] = 8'h00;
mem[16'hA129] = 8'hA1;
mem[16'hA12A] = 8'h00;
mem[16'hA12B] = 8'hA2;
mem[16'hA12C] = 8'h00;
mem[16'hA12D] = 8'h64;
mem[16'hA12E] = 8'h00;
mem[16'hA12F] = 8'h0A;
mem[16'hA130] = 8'h00;
mem[16'hA131] = 8'hA8;
mem[16'hA132] = 8'h00;
mem[16'hA133] = 8'h45;
mem[16'hA134] = 8'h00;
mem[16'hA135] = 8'h09;
mem[16'hA136] = 8'h00;
mem[16'hA137] = 8'h44;
mem[16'hA138] = 8'h00;
mem[16'hA139] = 8'h55;
mem[16'hA13A] = 8'h00;
mem[16'hA13B] = 8'h90;
mem[16'hA13C] = 8'h00;
mem[16'hA13D] = 8'hA5;
mem[16'hA13E] = 8'h00;
mem[16'hA13F] = 8'hD9;
mem[16'hA140] = 8'h00;
mem[16'hA141] = 8'hA9;
mem[16'hA142] = 8'h00;
mem[16'hA143] = 8'h0B;
mem[16'hA144] = 8'h00;
mem[16'hA145] = 8'h83;
mem[16'hA146] = 8'h00;
mem[16'hA147] = 8'h44;
mem[16'hA148] = 8'h00;
mem[16'hA149] = 8'h57;
mem[16'hA14A] = 8'h00;
mem[16'hA14B] = 8'h90;
mem[16'hA14C] = 8'h00;
mem[16'hA14D] = 8'hD0;
mem[16'hA14E] = 8'h00;
mem[16'hA14F] = 8'hAD;
mem[16'hA150] = 8'h00;
mem[16'hA151] = 8'hAA;
mem[16'hA152] = 8'h00;
mem[16'hA153] = 8'h94;
mem[16'hA154] = 8'h00;
mem[16'hA155] = 8'h4A;
mem[16'hA156] = 8'h00;
mem[16'hA157] = 8'hA5;
mem[16'hA158] = 8'h00;
mem[16'hA159] = 8'h99;
mem[16'hA15A] = 8'h00;
mem[16'hA15B] = 8'hAA;
mem[16'hA15C] = 8'h00;
mem[16'hA15D] = 8'h44;
mem[16'hA15E] = 8'h00;
mem[16'hA15F] = 8'h66;
mem[16'hA160] = 8'h00;
mem[16'hA161] = 8'h4C;
mem[16'hA162] = 8'h00;
mem[16'hA163] = 8'hA0;
mem[16'hA164] = 8'h00;
mem[16'hA165] = 8'hA9;
mem[16'hA166] = 8'h00;
mem[16'hA167] = 8'h0D;
mem[16'hA168] = 8'h00;
mem[16'hA169] = 8'hAA;
mem[16'hA16A] = 8'h00;
mem[16'hA16B] = 8'h65;
mem[16'hA16C] = 8'h00;
mem[16'hA16D] = 8'h68;
mem[16'hA16E] = 8'h00;
mem[16'hA16F] = 8'h7F;
mem[16'hA170] = 8'h00;
mem[16'hA171] = 8'h74;
mem[16'hA172] = 8'h00;
mem[16'hA173] = 8'h8D;
mem[16'hA174] = 8'h00;
mem[16'hA175] = 8'hAA;
mem[16'hA176] = 8'h00;
mem[16'hA177] = 8'hE9;
mem[16'hA178] = 8'h00;
mem[16'hA179] = 8'h9C;
mem[16'hA17A] = 8'h00;
mem[16'hA17B] = 8'h80;
mem[16'hA17C] = 8'h00;
mem[16'hA17D] = 8'h4C;
mem[16'hA17E] = 8'h00;
mem[16'hA17F] = 8'h9F;
mem[16'hA180] = 8'h00;
mem[16'hA181] = 8'h5B;
mem[16'hA182] = 8'h00;
mem[16'hA183] = 8'h20;
mem[16'hA184] = 8'h00;
mem[16'hA185] = 8'hA1;
mem[16'hA186] = 8'h00;
mem[16'hA187] = 8'h5F;
mem[16'hA188] = 8'h00;
mem[16'hA189] = 8'hAA;
mem[16'hA18A] = 8'h00;
mem[16'hA18B] = 8'h1F;
mem[16'hA18C] = 8'h00;
mem[16'hA18D] = 8'h48;
mem[16'hA18E] = 8'h00;
mem[16'hA18F] = 8'h1E;
mem[16'hA190] = 8'h00;
mem[16'hA191] = 8'h48;
mem[16'hA192] = 8'h00;
mem[16'hA193] = 8'hAE;
mem[16'hA194] = 8'h00;
mem[16'hA195] = 8'hAA;
mem[16'hA196] = 8'h00;
mem[16'hA197] = 8'h00;
mem[16'hA198] = 8'h00;
mem[16'hA199] = 8'hC9;
mem[16'hA19A] = 8'h00;
mem[16'hA19B] = 8'hF0;
mem[16'hA19C] = 8'h00;
mem[16'hA19D] = 8'hE8;
mem[16'hA19E] = 8'h00;
mem[16'hA19F] = 8'h5D;
mem[16'hA1A0] = 8'h00;
mem[16'hA1A1] = 8'hC9;
mem[16'hA1A2] = 8'h00;
mem[16'hA1A3] = 8'h60;
mem[16'hA1A4] = 8'h00;
mem[16'hA1A5] = 8'h93;
mem[16'hA1A6] = 8'h00;
mem[16'hA1A7] = 8'hF0;
mem[16'hA1A8] = 8'h00;
mem[16'hA1A9] = 8'hC9;
mem[16'hA1AA] = 8'h00;
mem[16'hA1AB] = 8'hF0;
mem[16'hA1AC] = 8'h00;
mem[16'hA1AD] = 8'h60;
mem[16'hA1AE] = 8'h00;
mem[16'hA1AF] = 8'h00;
mem[16'hA1B0] = 8'h00;
mem[16'hA1B1] = 8'h16;
mem[16'hA1B2] = 8'h00;
mem[16'hA1B3] = 8'hBA;
mem[16'hA1B4] = 8'h00;
mem[16'hA1B5] = 8'h88;
mem[16'hA1B6] = 8'h00;
mem[16'hA1B7] = 8'hFA;
mem[16'hA1B8] = 8'h00;
mem[16'hA1B9] = 8'hA9;
mem[16'hA1BA] = 8'h00;
mem[16'hA1BB] = 8'h85;
mem[16'hA1BC] = 8'h00;
mem[16'hA1BD] = 8'h85;
mem[16'hA1BE] = 8'h00;
mem[16'hA1BF] = 8'h20;
mem[16'hA1C0] = 8'h00;
mem[16'hA1C1] = 8'hA1;
mem[16'hA1C2] = 8'h00;
mem[16'hA1C3] = 8'hC9;
mem[16'hA1C4] = 8'h00;
mem[16'hA1C5] = 8'hF0;
mem[16'hA1C6] = 8'h00;
mem[16'hA1C7] = 8'h28;
mem[16'hA1C8] = 8'h00;
mem[16'hA1C9] = 8'hCE;
mem[16'hA1CA] = 8'h00;
mem[16'hA1CB] = 8'h20;
mem[16'hA1CC] = 8'h00;
mem[16'hA1CD] = 8'hA1;
mem[16'hA1CE] = 8'h00;
mem[16'hA1CF] = 8'h06;
mem[16'hA1D0] = 8'h00;
mem[16'hA1D1] = 8'h44;
mem[16'hA1D2] = 8'h00;
mem[16'hA1D3] = 8'h45;
mem[16'hA1D4] = 8'h00;
mem[16'hA1D5] = 8'h60;
mem[16'hA1D6] = 8'h00;
mem[16'hA1D7] = 8'hE9;
mem[16'hA1D8] = 8'h00;
mem[16'hA1D9] = 8'h30;
mem[16'hA1DA] = 8'h00;
mem[16'hA1DB] = 8'hC9;
mem[16'hA1DC] = 8'h00;
mem[16'hA1DD] = 8'hB0;
mem[16'hA1DE] = 8'h00;
mem[16'hA1DF] = 8'h20;
mem[16'hA1E0] = 8'h00;
mem[16'hA1E1] = 8'hA1;
mem[16'hA1E2] = 8'h00;
mem[16'hA1E3] = 8'h44;
mem[16'hA1E4] = 8'h00;
mem[16'hA1E5] = 8'hA9;
mem[16'hA1E6] = 8'h00;
mem[16'hA1E7] = 8'h65;
mem[16'hA1E8] = 8'h00;
mem[16'hA1E9] = 8'hA8;
mem[16'hA1EA] = 8'h00;
mem[16'hA1EB] = 8'hFE;
mem[16'hA1EC] = 8'h00;
mem[16'hA1ED] = 8'h20;
mem[16'hA1EE] = 8'h00;
mem[16'hA1EF] = 8'hA1;
mem[16'hA1F0] = 8'h00;
mem[16'hA1F1] = 8'h65;
mem[16'hA1F2] = 8'h00;
mem[16'hA1F3] = 8'h85;
mem[16'hA1F4] = 8'h00;
mem[16'hA1F5] = 8'h98;
mem[16'hA1F6] = 8'h00;
mem[16'hA1F7] = 8'h45;
mem[16'hA1F8] = 8'h00;
mem[16'hA1F9] = 8'h45;
mem[16'hA1FA] = 8'h00;
mem[16'hA1FB] = 8'hCF;
mem[16'hA1FC] = 8'h00;
mem[16'hA1FD] = 8'h60;
mem[16'hA1FE] = 8'h00;
mem[16'hA1FF] = 8'h44;
mem[16'hA200] = 8'h00;
mem[16'hA201] = 8'h45;
mem[16'hA202] = 8'h00;
mem[16'hA203] = 8'h28;
mem[16'hA204] = 8'h00;
mem[16'hA205] = 8'hA4;
mem[16'hA206] = 8'h00;
mem[16'hA207] = 8'hF0;
mem[16'hA208] = 8'h00;
mem[16'hA209] = 8'h38;
mem[16'hA20A] = 8'h00;
mem[16'hA20B] = 8'hB0;
mem[16'hA20C] = 8'h00;
mem[16'hA20D] = 8'hEE;
mem[16'hA20E] = 8'h00;
mem[16'hA20F] = 8'h0A;
mem[16'hA210] = 8'h00;
mem[16'hA211] = 8'h08;
mem[16'hA212] = 8'h00;
mem[16'hA213] = 8'h07;
mem[16'hA214] = 8'h00;
mem[16'hA215] = 8'hE6;
mem[16'hA216] = 8'h00;
mem[16'hA217] = 8'h10;
mem[16'hA218] = 8'h00;
mem[16'hA219] = 8'hE2;
mem[16'hA21A] = 8'h00;
mem[16'hA21B] = 8'h04;
mem[16'hA21C] = 8'h00;
mem[16'hA21D] = 8'hFE;
mem[16'hA21E] = 8'h00;
mem[16'hA21F] = 8'hCA;
mem[16'hA220] = 8'h00;
mem[16'hA221] = 8'hFA;
mem[16'hA222] = 8'h00;
mem[16'hA223] = 8'h44;
mem[16'hA224] = 8'h00;
mem[16'hA225] = 8'h44;
mem[16'hA226] = 8'h00;
mem[16'hA227] = 8'h04;
mem[16'hA228] = 8'h00;
mem[16'hA229] = 8'hA5;
mem[16'hA22A] = 8'h00;
mem[16'hA22B] = 8'h4C;
mem[16'hA22C] = 8'h00;
mem[16'hA22D] = 8'hFE;
mem[16'hA22E] = 8'h00;
mem[16'hA22F] = 8'h44;
mem[16'hA230] = 8'h00;
mem[16'hA231] = 8'h8B;
mem[16'hA232] = 8'h00;
mem[16'hA233] = 8'hAD;
mem[16'hA234] = 8'h00;
mem[16'hA235] = 8'hAA;
mem[16'hA236] = 8'h00;
mem[16'hA237] = 8'h74;
mem[16'hA238] = 8'h00;
mem[16'hA239] = 8'h8D;
mem[16'hA23A] = 8'h00;
mem[16'hA23B] = 8'hAA;
mem[16'hA23C] = 8'h00;
mem[16'hA23D] = 8'h2C;
mem[16'hA23E] = 8'h00;
mem[16'hA23F] = 8'hAA;
mem[16'hA240] = 8'h00;
mem[16'hA241] = 8'h03;
mem[16'hA242] = 8'h00;
mem[16'hA243] = 8'hC8;
mem[16'hA244] = 8'h00;
mem[16'hA245] = 8'hA9;
mem[16'hA246] = 8'h00;
mem[16'hA247] = 8'h4D;
mem[16'hA248] = 8'h00;
mem[16'hA249] = 8'hAA;
mem[16'hA24A] = 8'h00;
mem[16'hA24B] = 8'h5E;
mem[16'hA24C] = 8'h00;
mem[16'hA24D] = 8'h8D;
mem[16'hA24E] = 8'h00;
mem[16'hA24F] = 8'hAA;
mem[16'hA250] = 8'h00;
mem[16'hA251] = 8'hA9;
mem[16'hA252] = 8'h00;
mem[16'hA253] = 8'h8D;
mem[16'hA254] = 8'h00;
mem[16'hA255] = 8'hAA;
mem[16'hA256] = 8'h00;
mem[16'hA257] = 8'h44;
mem[16'hA258] = 8'h00;
mem[16'hA259] = 8'h20;
mem[16'hA25A] = 8'h00;
mem[16'hA25B] = 8'hA3;
mem[16'hA25C] = 8'h00;
mem[16'hA25D] = 8'h8D;
mem[16'hA25E] = 8'h00;
mem[16'hA25F] = 8'hAA;
mem[16'hA260] = 8'h00;
mem[16'hA261] = 8'hD4;
mem[16'hA262] = 8'h00;
mem[16'hA263] = 8'hA9;
mem[16'hA264] = 8'h00;
mem[16'hA265] = 8'h20;
mem[16'hA266] = 8'h00;
mem[16'hA267] = 8'hA2;
mem[16'hA268] = 8'h00;
mem[16'hA269] = 8'h64;
mem[16'hA26A] = 8'h00;
mem[16'hA26B] = 8'hA0;
mem[16'hA26C] = 8'h00;
mem[16'hA26D] = 8'h98;
mem[16'hA26E] = 8'h00;
mem[16'hA26F] = 8'h40;
mem[16'hA270] = 8'h00;
mem[16'hA271] = 8'hA9;
mem[16'hA272] = 8'h00;
mem[16'hA273] = 8'hD0;
mem[16'hA274] = 8'h00;
mem[16'hA275] = 8'hA9;
mem[16'hA276] = 8'h00;
mem[16'hA277] = 8'h20;
mem[16'hA278] = 8'h00;
mem[16'hA279] = 8'hA2;
mem[16'hA27A] = 8'h00;
mem[16'hA27B] = 8'hEA;
mem[16'hA27C] = 8'h00;
mem[16'hA27D] = 8'hA9;
mem[16'hA27E] = 8'h00;
mem[16'hA27F] = 8'hD0;
mem[16'hA280] = 8'h00;
mem[16'hA281] = 8'hAD;
mem[16'hA282] = 8'h00;
mem[16'hA283] = 8'h9D;
mem[16'hA284] = 8'h00;
mem[16'hA285] = 8'hBD;
mem[16'hA286] = 8'h00;
mem[16'hA287] = 8'hAD;
mem[16'hA288] = 8'h00;
mem[16'hA289] = 8'h9D;
mem[16'hA28A] = 8'h00;
mem[16'hA28B] = 8'hBE;
mem[16'hA28C] = 8'h00;
mem[16'hA28D] = 8'hA9;
mem[16'hA28E] = 8'h00;
mem[16'hA28F] = 8'h8D;
mem[16'hA290] = 8'h00;
mem[16'hA291] = 8'hAA;
mem[16'hA292] = 8'h00;
mem[16'hA293] = 8'hC8;
mem[16'hA294] = 8'h00;
mem[16'hA295] = 8'h4C;
mem[16'hA296] = 8'h00;
mem[16'hA297] = 8'hA2;
mem[16'hA298] = 8'h00;
mem[16'hA299] = 8'hA3;
mem[16'hA29A] = 8'h00;
mem[16'hA29B] = 8'h20;
mem[16'hA29C] = 8'h00;
mem[16'hA29D] = 8'hA6;
mem[16'hA29E] = 8'h00;
mem[16'hA29F] = 8'hFB;
mem[16'hA2A0] = 8'h00;
mem[16'hA2A1] = 8'h71;
mem[16'hA2A2] = 8'h00;
mem[16'hA2A3] = 8'hA9;
mem[16'hA2A4] = 8'h00;
mem[16'hA2A5] = 8'h4C;
mem[16'hA2A6] = 8'h00;
mem[16'hA2A7] = 8'hA3;
mem[16'hA2A8] = 8'h00;
mem[16'hA2A9] = 8'h01;
mem[16'hA2AA] = 8'h00;
mem[16'hA2AB] = 8'h63;
mem[16'hA2AC] = 8'h00;
mem[16'hA2AD] = 8'hAD;
mem[16'hA2AE] = 8'h00;
mem[16'hA2AF] = 8'hAA;
mem[16'hA2B0] = 8'h00;
mem[16'hA2B1] = 8'h0A;
mem[16'hA2B2] = 8'h00;
mem[16'hA2B3] = 8'h6D;
mem[16'hA2B4] = 8'h00;
mem[16'hA2B5] = 8'hD0;
mem[16'hA2B6] = 8'h00;
mem[16'hA2B7] = 8'hA9;
mem[16'hA2B8] = 8'h00;
mem[16'hA2B9] = 8'h8D;
mem[16'hA2BA] = 8'h00;
mem[16'hA2BB] = 8'hAA;
mem[16'hA2BC] = 8'h00;
mem[16'hA2BD] = 8'h6C;
mem[16'hA2BE] = 8'h00;
mem[16'hA2BF] = 8'h8D;
mem[16'hA2C0] = 8'h00;
mem[16'hA2C1] = 8'hB5;
mem[16'hA2C2] = 8'h00;
mem[16'hA2C3] = 8'h6D;
mem[16'hA2C4] = 8'h00;
mem[16'hA2C5] = 8'h8D;
mem[16'hA2C6] = 8'h00;
mem[16'hA2C7] = 8'hB5;
mem[16'hA2C8] = 8'h00;
mem[16'hA2C9] = 8'hEA;
mem[16'hA2CA] = 8'h00;
mem[16'hA2CB] = 8'hA5;
mem[16'hA2CC] = 8'h00;
mem[16'hA2CD] = 8'hD0;
mem[16'hA2CE] = 8'h00;
mem[16'hA2CF] = 8'h4C;
mem[16'hA2D0] = 8'h00;
mem[16'hA2D1] = 8'hA6;
mem[16'hA2D2] = 8'h00;
mem[16'hA2D3] = 8'h41;
mem[16'hA2D4] = 8'h00;
mem[16'hA2D5] = 8'h44;
mem[16'hA2D6] = 8'h00;
mem[16'hA2D7] = 8'h40;
mem[16'hA2D8] = 8'h00;
mem[16'hA2D9] = 8'h43;
mem[16'hA2DA] = 8'h00;
mem[16'hA2DB] = 8'h20;
mem[16'hA2DC] = 8'h00;
mem[16'hA2DD] = 8'hA7;
mem[16'hA2DE] = 8'h00;
mem[16'hA2DF] = 8'h1A;
mem[16'hA2E0] = 8'h00;
mem[16'hA2E1] = 8'hAD;
mem[16'hA2E2] = 8'h00;
mem[16'hA2E3] = 8'hAA;
mem[16'hA2E4] = 8'h00;
mem[16'hA2E5] = 8'hBB;
mem[16'hA2E6] = 8'h00;
mem[16'hA2E7] = 8'h4C;
mem[16'hA2E8] = 8'h00;
mem[16'hA2E9] = 8'hA6;
mem[16'hA2EA] = 8'h00;
mem[16'hA2EB] = 8'h75;
mem[16'hA2EC] = 8'h00;
mem[16'hA2ED] = 8'hC9;
mem[16'hA2EE] = 8'h00;
mem[16'hA2EF] = 8'hF0;
mem[16'hA2F0] = 8'h00;
mem[16'hA2F1] = 8'h20;
mem[16'hA2F2] = 8'h00;
mem[16'hA2F3] = 8'hA7;
mem[16'hA2F4] = 8'h00;
mem[16'hA2F5] = 8'h3A;
mem[16'hA2F6] = 8'h00;
mem[16'hA2F7] = 8'hFC;
mem[16'hA2F8] = 8'h00;
mem[16'hA2F9] = 8'h4C;
mem[16'hA2FA] = 8'h00;
mem[16'hA2FB] = 8'hA2;
mem[16'hA2FC] = 8'h00;
mem[16'hA2FD] = 8'hAF;
mem[16'hA2FE] = 8'h00;
mem[16'hA2FF] = 8'hD0;
mem[16'hA300] = 8'h00;
mem[16'hA301] = 8'hA9;
mem[16'hA302] = 8'h00;
mem[16'hA303] = 8'h8D;
mem[16'hA304] = 8'h00;
mem[16'hA305] = 8'hAA;
mem[16'hA306] = 8'h00;
mem[16'hA307] = 8'h00;
mem[16'hA308] = 8'h00;
mem[16'hA309] = 8'h91;
mem[16'hA30A] = 8'h00;
mem[16'hA30B] = 8'h20;
mem[16'hA30C] = 8'h00;
mem[16'hA30D] = 8'hA7;
mem[16'hA30E] = 8'h00;
mem[16'hA30F] = 8'h02;
mem[16'hA310] = 8'h00;
mem[16'hA311] = 8'hBB;
mem[16'hA312] = 8'h00;
mem[16'hA313] = 8'h4C;
mem[16'hA314] = 8'h00;
mem[16'hA315] = 8'hA6;
mem[16'hA316] = 8'h00;
mem[16'hA317] = 8'h92;
mem[16'hA318] = 8'h00;
mem[16'hA319] = 8'hD0;
mem[16'hA31A] = 8'h00;
mem[16'hA31B] = 8'h20;
mem[16'hA31C] = 8'h00;
mem[16'hA31D] = 8'hA7;
mem[16'hA31E] = 8'h00;
mem[16'hA31F] = 8'h10;
mem[16'hA320] = 8'h00;
mem[16'hA321] = 8'hAF;
mem[16'hA322] = 8'h00;
mem[16'hA323] = 8'hF0;
mem[16'hA324] = 8'h00;
mem[16'hA325] = 8'h20;
mem[16'hA326] = 8'h00;
mem[16'hA327] = 8'hA7;
mem[16'hA328] = 8'h00;
mem[16'hA329] = 8'hF1;
mem[16'hA32A] = 8'h00;
mem[16'hA32B] = 8'hFC;
mem[16'hA32C] = 8'h00;
mem[16'hA32D] = 8'h4C;
mem[16'hA32E] = 8'h00;
mem[16'hA32F] = 8'hA3;
mem[16'hA330] = 8'h00;
mem[16'hA331] = 8'hA9;
mem[16'hA332] = 8'h00;
mem[16'hA333] = 8'h2D;
mem[16'hA334] = 8'h00;
mem[16'hA335] = 8'hAA;
mem[16'hA336] = 8'h00;
mem[16'hA337] = 8'h09;
mem[16'hA338] = 8'h00;
mem[16'hA339] = 8'h03;
mem[16'hA33A] = 8'h00;
mem[16'hA33B] = 8'h00;
mem[16'hA33C] = 8'h00;
mem[16'hA33D] = 8'hA9;
mem[16'hA33E] = 8'h00;
mem[16'hA33F] = 8'h20;
mem[16'hA340] = 8'h00;
mem[16'hA341] = 8'hA3;
mem[16'hA342] = 8'h00;
mem[16'hA343] = 8'h73;
mem[16'hA344] = 8'h00;
mem[16'hA345] = 8'hAC;
mem[16'hA346] = 8'h00;
mem[16'hA347] = 8'hAA;
mem[16'hA348] = 8'h00;
mem[16'hA349] = 8'hE0;
mem[16'hA34A] = 8'h00;
mem[16'hA34B] = 8'hAD;
mem[16'hA34C] = 8'h00;
mem[16'hA34D] = 8'hAA;
mem[16'hA34E] = 8'h00;
mem[16'hA34F] = 8'h6C;
mem[16'hA350] = 8'h00;
mem[16'hA351] = 8'h20;
mem[16'hA352] = 8'h00;
mem[16'hA353] = 8'hA3;
mem[16'hA354] = 8'h00;
mem[16'hA355] = 8'h73;
mem[16'hA356] = 8'h00;
mem[16'hA357] = 8'hAC;
mem[16'hA358] = 8'h00;
mem[16'hA359] = 8'hAA;
mem[16'hA35A] = 8'h00;
mem[16'hA35B] = 8'hFF;
mem[16'hA35C] = 8'h00;
mem[16'hA35D] = 8'h20;
mem[16'hA35E] = 8'h00;
mem[16'hA35F] = 8'hA2;
mem[16'hA360] = 8'h00;
mem[16'hA361] = 8'h7F;
mem[16'hA362] = 8'h00;
mem[16'hA363] = 8'hC2;
mem[16'hA364] = 8'h00;
mem[16'hA365] = 8'hC9;
mem[16'hA366] = 8'h00;
mem[16'hA367] = 8'hF0;
mem[16'hA368] = 8'h00;
mem[16'hA369] = 8'h4C;
mem[16'hA36A] = 8'h00;
mem[16'hA36B] = 8'hA6;
mem[16'hA36C] = 8'h00;
mem[16'hA36D] = 8'h04;
mem[16'hA36E] = 8'h00;
mem[16'hA36F] = 8'hD5;
mem[16'hA370] = 8'h00;
mem[16'hA371] = 8'h20;
mem[16'hA372] = 8'h00;
mem[16'hA373] = 8'hA4;
mem[16'hA374] = 8'h00;
mem[16'hA375] = 8'hAD;
mem[16'hA376] = 8'h00;
mem[16'hA377] = 8'hAA;
mem[16'hA378] = 8'h00;
mem[16'hA379] = 8'h01;
mem[16'hA37A] = 8'h00;
mem[16'hA37B] = 8'h06;
mem[16'hA37C] = 8'h00;
mem[16'hA37D] = 8'h72;
mem[16'hA37E] = 8'h00;
mem[16'hA37F] = 8'h8C;
mem[16'hA380] = 8'h00;
mem[16'hA381] = 8'hAA;
mem[16'hA382] = 8'h00;
mem[16'hA383] = 8'h7A;
mem[16'hA384] = 8'h00;
mem[16'hA385] = 8'hAE;
mem[16'hA386] = 8'h00;
mem[16'hA387] = 8'hAA;
mem[16'hA388] = 8'h00;
mem[16'hA389] = 8'h73;
mem[16'hA38A] = 8'h00;
mem[16'hA38B] = 8'h4C;
mem[16'hA38C] = 8'h00;
mem[16'hA38D] = 8'hA4;
mem[16'hA38E] = 8'h00;
mem[16'hA38F] = 8'h5D;
mem[16'hA390] = 8'h00;
mem[16'hA391] = 8'h20;
mem[16'hA392] = 8'h00;
mem[16'hA393] = 8'hA8;
mem[16'hA394] = 8'h00;
mem[16'hA395] = 8'h72;
mem[16'hA396] = 8'h00;
mem[16'hA397] = 8'hAD;
mem[16'hA398] = 8'h00;
mem[16'hA399] = 8'hAA;
mem[16'hA39A] = 8'h00;
mem[16'hA39B] = 8'h20;
mem[16'hA39C] = 8'h00;
mem[16'hA39D] = 8'hD6;
mem[16'hA39E] = 8'h00;
mem[16'hA39F] = 8'h03;
mem[16'hA3A0] = 8'h00;
mem[16'hA3A1] = 8'hCC;
mem[16'hA3A2] = 8'h00;
mem[16'hA3A3] = 8'hA9;
mem[16'hA3A4] = 8'h00;
mem[16'hA3A5] = 8'h20;
mem[16'hA3A6] = 8'h00;
mem[16'hA3A7] = 8'hA3;
mem[16'hA3A8] = 8'h00;
mem[16'hA3A9] = 8'hA5;
mem[16'hA3AA] = 8'h00;
mem[16'hA3AB] = 8'hE5;
mem[16'hA3AC] = 8'h00;
mem[16'hA3AD] = 8'hA8;
mem[16'hA3AE] = 8'h00;
mem[16'hA3AF] = 8'hB0;
mem[16'hA3B0] = 8'h00;
mem[16'hA3B1] = 8'h68;
mem[16'hA3B2] = 8'h00;
mem[16'hA3B3] = 8'hE0;
mem[16'hA3B4] = 8'h00;
mem[16'hA3B5] = 8'hA5;
mem[16'hA3B6] = 8'h00;
mem[16'hA3B7] = 8'hA4;
mem[16'hA3B8] = 8'h00;
mem[16'hA3B9] = 8'h4C;
mem[16'hA3BA] = 8'h00;
mem[16'hA3BB] = 8'hA3;
mem[16'hA3BC] = 8'h00;
mem[16'hA3BD] = 8'h01;
mem[16'hA3BE] = 8'h00;
mem[16'hA3BF] = 8'hD5;
mem[16'hA3C0] = 8'h00;
mem[16'hA3C1] = 8'h38;
mem[16'hA3C2] = 8'h00;
mem[16'hA3C3] = 8'h4C;
mem[16'hA3C4] = 8'h00;
mem[16'hA3C5] = 8'hCA;
mem[16'hA3C6] = 8'h00;
mem[16'hA3C7] = 8'hA5;
mem[16'hA3C8] = 8'h00;
mem[16'hA3C9] = 8'hE5;
mem[16'hA3CA] = 8'h00;
mem[16'hA3CB] = 8'h20;
mem[16'hA3CC] = 8'h00;
mem[16'hA3CD] = 8'hA3;
mem[16'hA3CE] = 8'h00;
mem[16'hA3CF] = 8'hCB;
mem[16'hA3D0] = 8'h00;
mem[16'hA3D1] = 8'hCA;
mem[16'hA3D2] = 8'h00;
mem[16'hA3D3] = 8'hFF;
mem[16'hA3D4] = 8'h00;
mem[16'hA3D5] = 8'h8D;
mem[16'hA3D6] = 8'h00;
mem[16'hA3D7] = 8'hB5;
mem[16'hA3D8] = 8'h00;
mem[16'hA3D9] = 8'h20;
mem[16'hA3DA] = 8'h00;
mem[16'hA3DB] = 8'hA2;
mem[16'hA3DC] = 8'h00;
mem[16'hA3DD] = 8'h4C;
mem[16'hA3DE] = 8'h00;
mem[16'hA3DF] = 8'hA7;
mem[16'hA3E0] = 8'h00;
mem[16'hA3E1] = 8'hC1;
mem[16'hA3E2] = 8'h00;
mem[16'hA3E3] = 8'h8C;
mem[16'hA3E4] = 8'h00;
mem[16'hA3E5] = 8'hB5;
mem[16'hA3E6] = 8'h00;
mem[16'hA3E7] = 8'hC2;
mem[16'hA3E8] = 8'h00;
mem[16'hA3E9] = 8'hA9;
mem[16'hA3EA] = 8'h00;
mem[16'hA3EB] = 8'h8D;
mem[16'hA3EC] = 8'h00;
mem[16'hA3ED] = 8'hB5;
mem[16'hA3EE] = 8'h00;
mem[16'hA3EF] = 8'h01;
mem[16'hA3F0] = 8'h00;
mem[16'hA3F1] = 8'hBC;
mem[16'hA3F2] = 8'h00;
mem[16'hA3F3] = 8'h20;
mem[16'hA3F4] = 8'h00;
mem[16'hA3F5] = 8'hA6;
mem[16'hA3F6] = 8'h00;
mem[16'hA3F7] = 8'hC2;
mem[16'hA3F8] = 8'h00;
mem[16'hA3F9] = 8'h8D;
mem[16'hA3FA] = 8'h00;
mem[16'hA3FB] = 8'hB5;
mem[16'hA3FC] = 8'h00;
mem[16'hA3FD] = 8'hA8;
mem[16'hA3FE] = 8'h00;
mem[16'hA3FF] = 8'h8C;
mem[16'hA400] = 8'h00;
mem[16'hA401] = 8'hB5;
mem[16'hA402] = 8'h00;
mem[16'hA403] = 8'hC4;
mem[16'hA404] = 8'h00;
mem[16'hA405] = 8'hA9;
mem[16'hA406] = 8'h00;
mem[16'hA407] = 8'h4C;
mem[16'hA408] = 8'h00;
mem[16'hA409] = 8'hB6;
mem[16'hA40A] = 8'h00;
mem[16'hA40B] = 8'hA8;
mem[16'hA40C] = 8'h00;
mem[16'hA40D] = 8'h4C;
mem[16'hA40E] = 8'h00;
mem[16'hA40F] = 8'hA2;
mem[16'hA410] = 8'h00;
mem[16'hA411] = 8'hD0;
mem[16'hA412] = 8'h00;
mem[16'hA413] = 8'h20;
mem[16'hA414] = 8'h00;
mem[16'hA415] = 8'hA3;
mem[16'hA416] = 8'h00;
mem[16'hA417] = 8'hA8;
mem[16'hA418] = 8'h00;
mem[16'hA419] = 8'hA9;
mem[16'hA41A] = 8'h00;
mem[16'hA41B] = 8'h2D;
mem[16'hA41C] = 8'h00;
mem[16'hA41D] = 8'hB5;
mem[16'hA41E] = 8'h00;
mem[16'hA41F] = 8'hF0;
mem[16'hA420] = 8'h00;
mem[16'hA421] = 8'hC2;
mem[16'hA422] = 8'h00;
mem[16'hA423] = 8'hAD;
mem[16'hA424] = 8'h00;
mem[16'hA425] = 8'hAA;
mem[16'hA426] = 8'h00;
mem[16'hA427] = 8'h28;
mem[16'hA428] = 8'h00;
mem[16'hA429] = 8'h02;
mem[16'hA42A] = 8'h00;
mem[16'hA42B] = 8'hB1;
mem[16'hA42C] = 8'h00;
mem[16'hA42D] = 8'h20;
mem[16'hA42E] = 8'h00;
mem[16'hA42F] = 8'hA4;
mem[16'hA430] = 8'h00;
mem[16'hA431] = 8'h65;
mem[16'hA432] = 8'h00;
mem[16'hA433] = 8'hAA;
mem[16'hA434] = 8'h00;
mem[16'hA435] = 8'h65;
mem[16'hA436] = 8'h00;
mem[16'hA437] = 8'hC5;
mem[16'hA438] = 8'h00;
mem[16'hA439] = 8'hB0;
mem[16'hA43A] = 8'h00;
mem[16'hA43B] = 8'h85;
mem[16'hA43C] = 8'h00;
mem[16'hA43D] = 8'h85;
mem[16'hA43E] = 8'h00;
mem[16'hA43F] = 8'h86;
mem[16'hA440] = 8'h00;
mem[16'hA441] = 8'h86;
mem[16'hA442] = 8'h00;
mem[16'hA443] = 8'hA6;
mem[16'hA444] = 8'h00;
mem[16'hA445] = 8'hA4;
mem[16'hA446] = 8'h00;
mem[16'hA447] = 8'h20;
mem[16'hA448] = 8'h00;
mem[16'hA449] = 8'hA4;
mem[16'hA44A] = 8'h00;
mem[16'hA44B] = 8'h51;
mem[16'hA44C] = 8'h00;
mem[16'hA44D] = 8'h6C;
mem[16'hA44E] = 8'h00;
mem[16'hA44F] = 8'h9D;
mem[16'hA450] = 8'h00;
mem[16'hA451] = 8'h01;
mem[16'hA452] = 8'h00;
mem[16'hA453] = 8'hB1;
mem[16'hA454] = 8'h00;
mem[16'hA455] = 8'h20;
mem[16'hA456] = 8'h00;
mem[16'hA457] = 8'hA4;
mem[16'hA458] = 8'h00;
mem[16'hA459] = 8'hA5;
mem[16'hA45A] = 8'h00;
mem[16'hA45B] = 8'hED;
mem[16'hA45C] = 8'h00;
mem[16'hA45D] = 8'hAA;
mem[16'hA45E] = 8'h00;
mem[16'hA45F] = 8'hA5;
mem[16'hA460] = 8'h00;
mem[16'hA461] = 8'hED;
mem[16'hA462] = 8'h00;
mem[16'hA463] = 8'hAA;
mem[16'hA464] = 8'h00;
mem[16'hA465] = 8'h45;
mem[16'hA466] = 8'h00;
mem[16'hA467] = 8'hC4;
mem[16'hA468] = 8'h00;
mem[16'hA469] = 8'h90;
mem[16'hA46A] = 8'h00;
mem[16'hA46B] = 8'hF0;
mem[16'hA46C] = 8'h00;
mem[16'hA46D] = 8'h84;
mem[16'hA46E] = 8'h00;
mem[16'hA46F] = 8'h86;
mem[16'hA470] = 8'h00;
mem[16'hA471] = 8'h8E;
mem[16'hA472] = 8'h00;
mem[16'hA473] = 8'hB5;
mem[16'hA474] = 8'h00;
mem[16'hA475] = 8'hC4;
mem[16'hA476] = 8'h00;
mem[16'hA477] = 8'h4C;
mem[16'hA478] = 8'h00;
mem[16'hA479] = 8'hA4;
mem[16'hA47A] = 8'h00;
mem[16'hA47B] = 8'h0A;
mem[16'hA47C] = 8'h00;
mem[16'hA47D] = 8'h8D;
mem[16'hA47E] = 8'h00;
mem[16'hA47F] = 8'hB5;
mem[16'hA480] = 8'h00;
mem[16'hA481] = 8'h0B;
mem[16'hA482] = 8'h00;
mem[16'hA483] = 8'h8D;
mem[16'hA484] = 8'h00;
mem[16'hA485] = 8'hB5;
mem[16'hA486] = 8'h00;
mem[16'hA487] = 8'h00;
mem[16'hA488] = 8'h00;
mem[16'hA489] = 8'hC2;
mem[16'hA48A] = 8'h00;
mem[16'hA48B] = 8'hA9;
mem[16'hA48C] = 8'h00;
mem[16'hA48D] = 8'h8D;
mem[16'hA48E] = 8'h00;
mem[16'hA48F] = 8'hB5;
mem[16'hA490] = 8'h00;
mem[16'hA491] = 8'h03;
mem[16'hA492] = 8'h00;
mem[16'hA493] = 8'hBB;
mem[16'hA494] = 8'h00;
mem[16'hA495] = 8'hA9;
mem[16'hA496] = 8'h00;
mem[16'hA497] = 8'h8D;
mem[16'hA498] = 8'h00;
mem[16'hA499] = 8'hB5;
mem[16'hA49A] = 8'h00;
mem[16'hA49B] = 8'hA8;
mem[16'hA49C] = 8'h00;
mem[16'hA49D] = 8'hAD;
mem[16'hA49E] = 8'h00;
mem[16'hA49F] = 8'hAA;
mem[16'hA4A0] = 8'h00;
mem[16'hA4A1] = 8'hC2;
mem[16'hA4A2] = 8'h00;
mem[16'hA4A3] = 8'hA8;
mem[16'hA4A4] = 8'h00;
mem[16'hA4A5] = 8'h60;
mem[16'hA4A6] = 8'h00;
mem[16'hA4A7] = 8'h8D;
mem[16'hA4A8] = 8'h00;
mem[16'hA4A9] = 8'hB5;
mem[16'hA4AA] = 8'h00;
mem[16'hA4AB] = 8'h20;
mem[16'hA4AC] = 8'h00;
mem[16'hA4AD] = 8'hA2;
mem[16'hA4AE] = 8'h00;
mem[16'hA4AF] = 8'hCC;
mem[16'hA4B0] = 8'h00;
mem[16'hA4B1] = 8'hCD;
mem[16'hA4B2] = 8'h00;
mem[16'hA4B3] = 8'hB5;
mem[16'hA4B4] = 8'h00;
mem[16'hA4B5] = 8'h1A;
mem[16'hA4B6] = 8'h00;
mem[16'hA4B7] = 8'h5F;
mem[16'hA4B8] = 8'h00;
mem[16'hA4B9] = 8'h8E;
mem[16'hA4BA] = 8'h00;
mem[16'hA4BB] = 8'hAA;
mem[16'hA4BC] = 8'h00;
mem[16'hA4BD] = 8'hF0;
mem[16'hA4BE] = 8'h00;
mem[16'hA4BF] = 8'h4C;
mem[16'hA4C0] = 8'h00;
mem[16'hA4C1] = 8'hA5;
mem[16'hA4C2] = 8'h00;
mem[16'hA4C3] = 8'h1D;
mem[16'hA4C4] = 8'h00;
mem[16'hA4C5] = 8'h75;
mem[16'hA4C6] = 8'h00;
mem[16'hA4C7] = 8'h9D;
mem[16'hA4C8] = 8'h00;
mem[16'hA4C9] = 8'hAA;
mem[16'hA4CA] = 8'h00;
mem[16'hA4CB] = 8'h10;
mem[16'hA4CC] = 8'h00;
mem[16'hA4CD] = 8'h4C;
mem[16'hA4CE] = 8'h00;
mem[16'hA4CF] = 8'hA5;
mem[16'hA4D0] = 8'h00;
mem[16'hA4D1] = 8'hAD;
mem[16'hA4D2] = 8'h00;
mem[16'hA4D3] = 8'hAA;
mem[16'hA4D4] = 8'h00;
mem[16'hA4D5] = 8'h03;
mem[16'hA4D6] = 8'h00;
mem[16'hA4D7] = 8'hB7;
mem[16'hA4D8] = 8'h00;
mem[16'hA4D9] = 8'h20;
mem[16'hA4DA] = 8'h00;
mem[16'hA4DB] = 8'hA4;
mem[16'hA4DC] = 8'h00;
mem[16'hA4DD] = 8'hC8;
mem[16'hA4DE] = 8'h00;
mem[16'hA4DF] = 8'h20;
mem[16'hA4E0] = 8'h00;
mem[16'hA4E1] = 8'hA8;
mem[16'hA4E2] = 8'h00;
mem[16'hA4E3] = 8'h58;
mem[16'hA4E4] = 8'h00;
mem[16'hA4E5] = 8'hA5;
mem[16'hA4E6] = 8'h00;
mem[16'hA4E7] = 8'h85;
mem[16'hA4E8] = 8'h00;
mem[16'hA4E9] = 8'hA5;
mem[16'hA4EA] = 8'h00;
mem[16'hA4EB] = 8'h85;
mem[16'hA4EC] = 8'h00;
mem[16'hA4ED] = 8'h6C;
mem[16'hA4EE] = 8'h00;
mem[16'hA4EF] = 8'h9D;
mem[16'hA4F0] = 8'h00;
mem[16'hA4F1] = 8'h16;
mem[16'hA4F2] = 8'h00;
mem[16'hA4F3] = 8'h20;
mem[16'hA4F4] = 8'h00;
mem[16'hA4F5] = 8'h9F;
mem[16'hA4F6] = 8'h00;
mem[16'hA4F7] = 8'h51;
mem[16'hA4F8] = 8'h00;
mem[16'hA4F9] = 8'h6C;
mem[16'hA4FA] = 8'h00;
mem[16'hA4FB] = 8'h9D;
mem[16'hA4FC] = 8'h00;
mem[16'hA4FD] = 8'h65;
mem[16'hA4FE] = 8'h00;
mem[16'hA4FF] = 8'h85;
mem[16'hA500] = 8'h00;
mem[16'hA501] = 8'h85;
mem[16'hA502] = 8'h00;
mem[16'hA503] = 8'h4C;
mem[16'hA504] = 8'h00;
mem[16'hA505] = 8'hD7;
mem[16'hA506] = 8'h00;
mem[16'hA507] = 8'h65;
mem[16'hA508] = 8'h00;
mem[16'hA509] = 8'h85;
mem[16'hA50A] = 8'h00;
mem[16'hA50B] = 8'h85;
mem[16'hA50C] = 8'h00;
mem[16'hA50D] = 8'h4C;
mem[16'hA50E] = 8'h00;
mem[16'hA50F] = 8'h0F;
mem[16'hA510] = 8'h00;
mem[16'hA511] = 8'h26;
mem[16'hA512] = 8'h00;
mem[16'hA513] = 8'hA9;
mem[16'hA514] = 8'h00;
mem[16'hA515] = 8'h8D;
mem[16'hA516] = 8'h00;
mem[16'hA517] = 8'hAA;
mem[16'hA518] = 8'h00;
mem[16'hA519] = 8'h83;
mem[16'hA51A] = 8'h00;
mem[16'hA51B] = 8'h20;
mem[16'hA51C] = 8'h00;
mem[16'hA51D] = 8'hA5;
mem[16'hA51E] = 8'h00;
mem[16'hA51F] = 8'h01;
mem[16'hA520] = 8'h00;
mem[16'hA521] = 8'h51;
mem[16'hA522] = 8'h00;
mem[16'hA523] = 8'h4C;
mem[16'hA524] = 8'h00;
mem[16'hA525] = 8'h9F;
mem[16'hA526] = 8'h00;
mem[16'hA527] = 8'h64;
mem[16'hA528] = 8'h00;
mem[16'hA529] = 8'h90;
mem[16'hA52A] = 8'h00;
mem[16'hA52B] = 8'h20;
mem[16'hA52C] = 8'h00;
mem[16'hA52D] = 8'hA2;
mem[16'hA52E] = 8'h00;
mem[16'hA52F] = 8'h34;
mem[16'hA530] = 8'h00;
mem[16'hA531] = 8'h20;
mem[16'hA532] = 8'h00;
mem[16'hA533] = 8'hA7;
mem[16'hA534] = 8'h00;
mem[16'hA535] = 8'h65;
mem[16'hA536] = 8'h00;
mem[16'hA537] = 8'h29;
mem[16'hA538] = 8'h00;
mem[16'hA539] = 8'hF0;
mem[16'hA53A] = 8'h00;
mem[16'hA53B] = 8'hA2;
mem[16'hA53C] = 8'h00;
mem[16'hA53D] = 8'hBD;
mem[16'hA53E] = 8'h00;
mem[16'hA53F] = 8'hAA;
mem[16'hA540] = 8'h00;
mem[16'hA541] = 8'hBD;
mem[16'hA542] = 8'h00;
mem[16'hA543] = 8'hCA;
mem[16'hA544] = 8'h00;
mem[16'hA545] = 8'hF7;
mem[16'hA546] = 8'h00;
mem[16'hA547] = 8'h0A;
mem[16'hA548] = 8'h00;
mem[16'hA549] = 8'hBB;
mem[16'hA54A] = 8'h00;
mem[16'hA54B] = 8'h20;
mem[16'hA54C] = 8'h00;
mem[16'hA54D] = 8'hA6;
mem[16'hA54E] = 8'h00;
mem[16'hA54F] = 8'hA9;
mem[16'hA550] = 8'h00;
mem[16'hA551] = 8'h2D;
mem[16'hA552] = 8'h00;
mem[16'hA553] = 8'hAA;
mem[16'hA554] = 8'h00;
mem[16'hA555] = 8'h05;
mem[16'hA556] = 8'h00;
mem[16'hA557] = 8'h66;
mem[16'hA558] = 8'h00;
mem[16'hA559] = 8'hD0;
mem[16'hA55A] = 8'h00;
mem[16'hA55B] = 8'hA9;
mem[16'hA55C] = 8'h00;
mem[16'hA55D] = 8'h8D;
mem[16'hA55E] = 8'h00;
mem[16'hA55F] = 8'hAA;
mem[16'hA560] = 8'h00;
mem[16'hA561] = 8'h0D;
mem[16'hA562] = 8'h00;
mem[16'hA563] = 8'h8D;
mem[16'hA564] = 8'h00;
mem[16'hA565] = 8'hB5;
mem[16'hA566] = 8'h00;
mem[16'hA567] = 8'h0B;
mem[16'hA568] = 8'h00;
mem[16'hA569] = 8'hAA;
mem[16'hA56A] = 8'h00;
mem[16'hA56B] = 8'h4C;
mem[16'hA56C] = 8'h00;
mem[16'hA56D] = 8'hA3;
mem[16'hA56E] = 8'h00;
mem[16'hA56F] = 8'h06;
mem[16'hA570] = 8'h00;
mem[16'hA571] = 8'hAA;
mem[16'hA572] = 8'h00;
mem[16'hA573] = 8'hAD;
mem[16'hA574] = 8'h00;
mem[16'hA575] = 8'hB5;
mem[16'hA576] = 8'h00;
mem[16'hA577] = 8'h66;
mem[16'hA578] = 8'h00;
mem[16'hA579] = 8'h60;
mem[16'hA57A] = 8'h00;
mem[16'hA57B] = 8'h4C;
mem[16'hA57C] = 8'h00;
mem[16'hA57D] = 8'hB2;
mem[16'hA57E] = 8'h00;
mem[16'hA57F] = 8'hF0;
mem[16'hA580] = 8'h00;
mem[16'hA581] = 8'hA9;
mem[16'hA582] = 8'h00;
mem[16'hA583] = 8'h8D;
mem[16'hA584] = 8'h00;
mem[16'hA585] = 8'hAA;
mem[16'hA586] = 8'h00;
mem[16'hA587] = 8'h1E;
mem[16'hA588] = 8'h00;
mem[16'hA589] = 8'h97;
mem[16'hA58A] = 8'h00;
mem[16'hA58B] = 8'hA2;
mem[16'hA58C] = 8'h00;
mem[16'hA58D] = 8'hBD;
mem[16'hA58E] = 8'h00;
mem[16'hA58F] = 8'hAA;
mem[16'hA590] = 8'h00;
mem[16'hA591] = 8'h74;
mem[16'hA592] = 8'h00;
mem[16'hA593] = 8'hCA;
mem[16'hA594] = 8'h00;
mem[16'hA595] = 8'hF7;
mem[16'hA596] = 8'h00;
mem[16'hA597] = 8'hC0;
mem[16'hA598] = 8'h00;
mem[16'hA599] = 8'h51;
mem[16'hA59A] = 8'h00;
mem[16'hA59B] = 8'h4C;
mem[16'hA59C] = 8'h00;
mem[16'hA59D] = 8'hA4;
mem[16'hA59E] = 8'h00;
mem[16'hA59F] = 8'h20;
mem[16'hA5A0] = 8'h00;
mem[16'hA5A1] = 8'hB2;
mem[16'hA5A2] = 8'h00;
mem[16'hA5A3] = 8'hF0;
mem[16'hA5A4] = 8'h00;
mem[16'hA5A5] = 8'hA9;
mem[16'hA5A6] = 8'h00;
mem[16'hA5A7] = 8'h4C;
mem[16'hA5A8] = 8'h00;
mem[16'hA5A9] = 8'hA6;
mem[16'hA5AA] = 8'h00;
mem[16'hA5AB] = 8'h00;
mem[16'hA5AC] = 8'h00;
mem[16'hA5AD] = 8'hB7;
mem[16'hA5AE] = 8'h00;
mem[16'hA5AF] = 8'h4C;
mem[16'hA5B0] = 8'h00;
mem[16'hA5B1] = 8'h9D;
mem[16'hA5B2] = 8'h00;
mem[16'hA5B3] = 8'h00;
mem[16'hA5B4] = 8'h00;
mem[16'hA5B5] = 8'hF0;
mem[16'hA5B6] = 8'h00;
mem[16'hA5B7] = 8'h8D;
mem[16'hA5B8] = 8'h00;
mem[16'hA5B9] = 8'hC0;
mem[16'hA5BA] = 8'h00;
mem[16'hA5BB] = 8'h00;
mem[16'hA5BC] = 8'h00;
mem[16'hA5BD] = 8'hF0;
mem[16'hA5BE] = 8'h00;
mem[16'hA5BF] = 8'h8D;
mem[16'hA5C0] = 8'h00;
mem[16'hA5C1] = 8'hC0;
mem[16'hA5C2] = 8'h00;
mem[16'hA5C3] = 8'h00;
mem[16'hA5C4] = 8'h00;
mem[16'hA5C5] = 8'h60;
mem[16'hA5C6] = 8'h00;
mem[16'hA5C7] = 8'hA3;
mem[16'hA5C8] = 8'h00;
mem[16'hA5C9] = 8'hAD;
mem[16'hA5CA] = 8'h00;
mem[16'hA5CB] = 8'hAA;
mem[16'hA5CC] = 8'h00;
mem[16'hA5CD] = 8'hB4;
mem[16'hA5CE] = 8'h00;
mem[16'hA5CF] = 8'hAD;
mem[16'hA5D0] = 8'h00;
mem[16'hA5D1] = 8'hAA;
mem[16'hA5D2] = 8'h00;
mem[16'hA5D3] = 8'hB5;
mem[16'hA5D4] = 8'h00;
mem[16'hA5D5] = 8'hAD;
mem[16'hA5D6] = 8'h00;
mem[16'hA5D7] = 8'hAA;
mem[16'hA5D8] = 8'h00;
mem[16'hA5D9] = 8'hB3;
mem[16'hA5DA] = 8'h00;
mem[16'hA5DB] = 8'hD0;
mem[16'hA5DC] = 8'h00;
mem[16'hA5DD] = 8'h20;
mem[16'hA5DE] = 8'h00;
mem[16'hA5DF] = 8'hA7;
mem[16'hA5E0] = 8'h00;
mem[16'hA5E1] = 8'h06;
mem[16'hA5E2] = 8'h00;
mem[16'hA5E3] = 8'hA3;
mem[16'hA5E4] = 8'h00;
mem[16'hA5E5] = 8'h4C;
mem[16'hA5E6] = 8'h00;
mem[16'hA5E7] = 8'hA5;
mem[16'hA5E8] = 8'h00;
mem[16'hA5E9] = 8'h4E;
mem[16'hA5EA] = 8'h00;
mem[16'hA5EB] = 8'hAD;
mem[16'hA5EC] = 8'h00;
mem[16'hA5ED] = 8'hAA;
mem[16'hA5EE] = 8'h00;
mem[16'hA5EF] = 8'h04;
mem[16'hA5F0] = 8'h00;
mem[16'hA5F1] = 8'h1B;
mem[16'hA5F2] = 8'h00;
mem[16'hA5F3] = 8'h6E;
mem[16'hA5F4] = 8'h00;
mem[16'hA5F5] = 8'hD0;
mem[16'hA5F6] = 8'h00;
mem[16'hA5F7] = 8'hAE;
mem[16'hA5F8] = 8'h00;
mem[16'hA5F9] = 8'hAA;
mem[16'hA5FA] = 8'h00;
mem[16'hA5FB] = 8'h11;
mem[16'hA5FC] = 8'h00;
mem[16'hA5FD] = 8'h6F;
mem[16'hA5FE] = 8'h00;
mem[16'hA5FF] = 8'hCE;
mem[16'hA600] = 8'h00;
mem[16'hA601] = 8'hAA;
mem[16'hA602] = 8'h00;
mem[16'hA603] = 8'h8C;
mem[16'hA604] = 8'h00;
mem[16'hA605] = 8'hF0;
mem[16'hA606] = 8'h00;
mem[16'hA607] = 8'hC9;
mem[16'hA608] = 8'h00;
mem[16'hA609] = 8'hD0;
mem[16'hA60A] = 8'h00;
mem[16'hA60B] = 8'hF0;
mem[16'hA60C] = 8'h00;
mem[16'hA60D] = 8'h60;
mem[16'hA60E] = 8'h00;
mem[16'hA60F] = 8'h5E;
mem[16'hA610] = 8'h00;
mem[16'hA611] = 8'hB0;
mem[16'hA612] = 8'h00;
mem[16'hA613] = 8'hAD;
mem[16'hA614] = 8'h00;
mem[16'hA615] = 8'hAA;
mem[16'hA616] = 8'h00;
mem[16'hA617] = 8'hC3;
mem[16'hA618] = 8'h00;
mem[16'hA619] = 8'hA9;
mem[16'hA61A] = 8'h00;
mem[16'hA61B] = 8'h8D;
mem[16'hA61C] = 8'h00;
mem[16'hA61D] = 8'hB5;
mem[16'hA61E] = 8'h00;
mem[16'hA61F] = 8'h01;
mem[16'hA620] = 8'h00;
mem[16'hA621] = 8'hBC;
mem[16'hA622] = 8'h00;
mem[16'hA623] = 8'h4C;
mem[16'hA624] = 8'h00;
mem[16'hA625] = 8'hA6;
mem[16'hA626] = 8'h00;
mem[16'hA627] = 8'h5E;
mem[16'hA628] = 8'h00;
mem[16'hA629] = 8'hB0;
mem[16'hA62A] = 8'h00;
mem[16'hA62B] = 8'hA9;
mem[16'hA62C] = 8'h00;
mem[16'hA62D] = 8'h8D;
mem[16'hA62E] = 8'h00;
mem[16'hA62F] = 8'hAA;
mem[16'hA630] = 8'h00;
mem[16'hA631] = 8'h8C;
mem[16'hA632] = 8'h00;
mem[16'hA633] = 8'hD0;
mem[16'hA634] = 8'h00;
mem[16'hA635] = 8'h20;
mem[16'hA636] = 8'h00;
mem[16'hA637] = 8'hA2;
mem[16'hA638] = 8'h00;
mem[16'hA639] = 8'h03;
mem[16'hA63A] = 8'h00;
mem[16'hA63B] = 8'h52;
mem[16'hA63C] = 8'h00;
mem[16'hA63D] = 8'hF0;
mem[16'hA63E] = 8'h00;
mem[16'hA63F] = 8'hA9;
mem[16'hA640] = 8'h00;
mem[16'hA641] = 8'h4C;
mem[16'hA642] = 8'h00;
mem[16'hA643] = 8'hA6;
mem[16'hA644] = 8'h00;
mem[16'hA645] = 8'hE0;
mem[16'hA646] = 8'h00;
mem[16'hA647] = 8'h02;
mem[16'hA648] = 8'h00;
mem[16'hA649] = 8'h7F;
mem[16'hA64A] = 8'h00;
mem[16'hA64B] = 8'h5C;
mem[16'hA64C] = 8'h00;
mem[16'hA64D] = 8'hAE;
mem[16'hA64E] = 8'h00;
mem[16'hA64F] = 8'hAA;
mem[16'hA650] = 8'h00;
mem[16'hA651] = 8'h09;
mem[16'hA652] = 8'h00;
mem[16'hA653] = 8'hBD;
mem[16'hA654] = 8'h00;
mem[16'hA655] = 8'h02;
mem[16'hA656] = 8'h00;
mem[16'hA657] = 8'h80;
mem[16'hA658] = 8'h00;
mem[16'hA659] = 8'h00;
mem[16'hA65A] = 8'h00;
mem[16'hA65B] = 8'h4C;
mem[16'hA65C] = 8'h00;
mem[16'hA65D] = 8'h9F;
mem[16'hA65E] = 8'h00;
mem[16'hA65F] = 8'hAD;
mem[16'hA660] = 8'h00;
mem[16'hA661] = 8'hAA;
mem[16'hA662] = 8'h00;
mem[16'hA663] = 8'h0E;
mem[16'hA664] = 8'h00;
mem[16'hA665] = 8'h76;
mem[16'hA666] = 8'h00;
mem[16'hA667] = 8'hF0;
mem[16'hA668] = 8'h00;
mem[16'hA669] = 8'hA6;
mem[16'hA66A] = 8'h00;
mem[16'hA66B] = 8'hE0;
mem[16'hA66C] = 8'h00;
mem[16'hA66D] = 8'hF0;
mem[16'hA66E] = 8'h00;
mem[16'hA66F] = 8'h68;
mem[16'hA670] = 8'h00;
mem[16'hA671] = 8'h60;
mem[16'hA672] = 8'h00;
mem[16'hA673] = 8'hD9;
mem[16'hA674] = 8'h00;
mem[16'hA675] = 8'hF9;
mem[16'hA676] = 8'h00;
mem[16'hA677] = 8'h38;
mem[16'hA678] = 8'h00;
mem[16'hA679] = 8'h20;
mem[16'hA67A] = 8'h00;
mem[16'hA67B] = 8'hA2;
mem[16'hA67C] = 8'h00;
mem[16'hA67D] = 8'h5B;
mem[16'hA67E] = 8'h00;
mem[16'hA67F] = 8'h4C;
mem[16'hA680] = 8'h00;
mem[16'hA681] = 8'h9F;
mem[16'hA682] = 8'h00;
mem[16'hA683] = 8'h9D;
mem[16'hA684] = 8'h00;
mem[16'hA685] = 8'h20;
mem[16'hA686] = 8'h00;
mem[16'hA687] = 8'hA7;
mem[16'hA688] = 8'h00;
mem[16'hA689] = 8'h03;
mem[16'hA68A] = 8'h00;
mem[16'hA68B] = 8'hA1;
mem[16'hA68C] = 8'h00;
mem[16'hA68D] = 8'h03;
mem[16'hA68E] = 8'h00;
mem[16'hA68F] = 8'hBB;
mem[16'hA690] = 8'h00;
mem[16'hA691] = 8'hA9;
mem[16'hA692] = 8'h00;
mem[16'hA693] = 8'h8D;
mem[16'hA694] = 8'h00;
mem[16'hA695] = 8'hB5;
mem[16'hA696] = 8'h00;
mem[16'hA697] = 8'hA8;
mem[16'hA698] = 8'h00;
mem[16'hA699] = 8'hAD;
mem[16'hA69A] = 8'h00;
mem[16'hA69B] = 8'hB5;
mem[16'hA69C] = 8'h00;
mem[16'hA69D] = 8'hAD;
mem[16'hA69E] = 8'h00;
mem[16'hA69F] = 8'hAA;
mem[16'hA6A0] = 8'h00;
mem[16'hA6A1] = 8'h41;
mem[16'hA6A2] = 8'h00;
mem[16'hA6A3] = 8'hB4;
mem[16'hA6A4] = 8'h00;
mem[16'hA6A5] = 8'h85;
mem[16'hA6A6] = 8'h00;
mem[16'hA6A7] = 8'h60;
mem[16'hA6A8] = 8'h00;
mem[16'hA6A9] = 8'h06;
mem[16'hA6AA] = 8'h00;
mem[16'hA6AB] = 8'h90;
mem[16'hA6AC] = 8'h00;
mem[16'hA6AD] = 8'hAD;
mem[16'hA6AE] = 8'h00;
mem[16'hA6AF] = 8'hB5;
mem[16'hA6B0] = 8'h00;
mem[16'hA6B1] = 8'h05;
mem[16'hA6B2] = 8'h00;
mem[16'hA6B3] = 8'h03;
mem[16'hA6B4] = 8'h00;
mem[16'hA6B5] = 8'h5E;
mem[16'hA6B6] = 8'h00;
mem[16'hA6B7] = 8'h4C;
mem[16'hA6B8] = 8'h00;
mem[16'hA6B9] = 8'hB6;
mem[16'hA6BA] = 8'h00;
mem[16'hA6BB] = 8'hEA;
mem[16'hA6BC] = 8'h00;
mem[16'hA6BD] = 8'hEA;
mem[16'hA6BE] = 8'h00;
mem[16'hA6BF] = 8'h00;
mem[16'hA6C0] = 8'h00;
mem[16'hA6C1] = 8'hC3;
mem[16'hA6C2] = 8'h00;
mem[16'hA6C3] = 8'h60;
mem[16'hA6C4] = 8'h00;
mem[16'hA6C5] = 8'h0B;
mem[16'hA6C6] = 8'h00;
mem[16'hA6C7] = 8'h0A;
mem[16'hA6C8] = 8'h00;
mem[16'hA6C9] = 8'h0C;
mem[16'hA6CA] = 8'h00;
mem[16'hA6CB] = 8'h06;
mem[16'hA6CC] = 8'h00;
mem[16'hA6CD] = 8'h0E;
mem[16'hA6CE] = 8'h00;
mem[16'hA6CF] = 8'h02;
mem[16'hA6D0] = 8'h00;
mem[16'hA6D1] = 8'h0D;
mem[16'hA6D2] = 8'h00;
mem[16'hA6D3] = 8'h5C;
mem[16'hA6D4] = 8'h00;
mem[16'hA6D5] = 8'h20;
mem[16'hA6D6] = 8'h00;
mem[16'hA6D7] = 8'hBF;
mem[16'hA6D8] = 8'h00;
mem[16'hA6D9] = 8'hB6;
mem[16'hA6DA] = 8'h00;
mem[16'hA6DB] = 8'hF0;
mem[16'hA6DC] = 8'h00;
mem[16'hA6DD] = 8'hA5;
mem[16'hA6DE] = 8'h00;
mem[16'hA6DF] = 8'h30;
mem[16'hA6E0] = 8'h00;
mem[16'hA6E1] = 8'hA2;
mem[16'hA6E2] = 8'h00;
mem[16'hA6E3] = 8'h20;
mem[16'hA6E4] = 8'h00;
mem[16'hA6E5] = 8'hA7;
mem[16'hA6E6] = 8'h00;
mem[16'hA6E7] = 8'h5C;
mem[16'hA6E8] = 8'h00;
mem[16'hA6E9] = 8'h20;
mem[16'hA6EA] = 8'h00;
mem[16'hA6EB] = 8'hA7;
mem[16'hA6EC] = 8'h00;
mem[16'hA6ED] = 8'hC8;
mem[16'hA6EE] = 8'h00;
mem[16'hA6EF] = 8'h20;
mem[16'hA6F0] = 8'h00;
mem[16'hA6F1] = 8'hA8;
mem[16'hA6F2] = 8'h00;
mem[16'hA6F3] = 8'h5E;
mem[16'hA6F4] = 8'h00;
mem[16'hA6F5] = 8'hAE;
mem[16'hA6F6] = 8'h00;
mem[16'hA6F7] = 8'hAA;
mem[16'hA6F8] = 8'h00;
mem[16'hA6F9] = 8'h03;
mem[16'hA6FA] = 8'h00;
mem[16'hA6FB] = 8'h03;
mem[16'hA6FC] = 8'h00;
mem[16'hA6FD] = 8'h5A;
mem[16'hA6FE] = 8'h00;
mem[16'hA6FF] = 8'h6C;
mem[16'hA700] = 8'h00;
mem[16'hA701] = 8'h9D;
mem[16'hA702] = 8'h00;
mem[16'hA703] = 8'h3F;
mem[16'hA704] = 8'h00;
mem[16'hA705] = 8'hAA;
mem[16'hA706] = 8'h00;
mem[16'hA707] = 8'h63;
mem[16'hA708] = 8'h00;
mem[16'hA709] = 8'hBD;
mem[16'hA70A] = 8'h00;
mem[16'hA70B] = 8'hA9;
mem[16'hA70C] = 8'h00;
mem[16'hA70D] = 8'h09;
mem[16'hA70E] = 8'h00;
mem[16'hA70F] = 8'h20;
mem[16'hA710] = 8'h00;
mem[16'hA711] = 8'h9F;
mem[16'hA712] = 8'h00;
mem[16'hA713] = 8'h63;
mem[16'hA714] = 8'h00;
mem[16'hA715] = 8'hE8;
mem[16'hA716] = 8'h00;
mem[16'hA717] = 8'h10;
mem[16'hA718] = 8'h00;
mem[16'hA719] = 8'h60;
mem[16'hA71A] = 8'h00;
mem[16'hA71B] = 8'h66;
mem[16'hA71C] = 8'h00;
mem[16'hA71D] = 8'h8D;
mem[16'hA71E] = 8'h00;
mem[16'hA71F] = 8'hB5;
mem[16'hA720] = 8'h00;
mem[16'hA721] = 8'h68;
mem[16'hA722] = 8'h00;
mem[16'hA723] = 8'h8D;
mem[16'hA724] = 8'h00;
mem[16'hA725] = 8'hB5;
mem[16'hA726] = 8'h00;
mem[16'hA727] = 8'h6A;
mem[16'hA728] = 8'h00;
mem[16'hA729] = 8'h8D;
mem[16'hA72A] = 8'h00;
mem[16'hA72B] = 8'hB5;
mem[16'hA72C] = 8'h00;
mem[16'hA72D] = 8'h06;
mem[16'hA72E] = 8'h00;
mem[16'hA72F] = 8'h8D;
mem[16'hA730] = 8'h00;
mem[16'hA731] = 8'hB5;
mem[16'hA732] = 8'h00;
mem[16'hA733] = 8'h07;
mem[16'hA734] = 8'h00;
mem[16'hA735] = 8'h8D;
mem[16'hA736] = 8'h00;
mem[16'hA737] = 8'hB5;
mem[16'hA738] = 8'h00;
mem[16'hA739] = 8'h40;
mem[16'hA73A] = 8'h00;
mem[16'hA73B] = 8'h4F;
mem[16'hA73C] = 8'h00;
mem[16'hA73D] = 8'hA5;
mem[16'hA73E] = 8'h00;
mem[16'hA73F] = 8'h8D;
mem[16'hA740] = 8'h00;
mem[16'hA741] = 8'hAA;
mem[16'hA742] = 8'h00;
mem[16'hA743] = 8'hA0;
mem[16'hA744] = 8'h00;
mem[16'hA745] = 8'hB9;
mem[16'hA746] = 8'h00;
mem[16'hA747] = 8'hAA;
mem[16'hA748] = 8'h00;
mem[16'hA749] = 8'h40;
mem[16'hA74A] = 8'h00;
mem[16'hA74B] = 8'h10;
mem[16'hA74C] = 8'h00;
mem[16'hA74D] = 8'h60;
mem[16'hA74E] = 8'h00;
mem[16'hA74F] = 8'h1E;
mem[16'hA750] = 8'h00;
mem[16'hA751] = 8'h40;
mem[16'hA752] = 8'h00;
mem[16'hA753] = 8'hA9;
mem[16'hA754] = 8'h00;
mem[16'hA755] = 8'hC8;
mem[16'hA756] = 8'h00;
mem[16'hA757] = 8'h26;
mem[16'hA758] = 8'h00;
mem[16'hA759] = 8'hF6;
mem[16'hA75A] = 8'h00;
mem[16'hA75B] = 8'hA0;
mem[16'hA75C] = 8'h00;
mem[16'hA75D] = 8'h8C;
mem[16'hA75E] = 8'h00;
mem[16'hA75F] = 8'hAA;
mem[16'hA760] = 8'h00;
mem[16'hA761] = 8'h52;
mem[16'hA762] = 8'h00;
mem[16'hA763] = 8'h60;
mem[16'hA764] = 8'h00;
mem[16'hA765] = 8'h00;
mem[16'hA766] = 8'h00;
mem[16'hA767] = 8'h45;
mem[16'hA768] = 8'h00;
mem[16'hA769] = 8'h92;
mem[16'hA76A] = 8'h00;
mem[16'hA76B] = 8'h4C;
mem[16'hA76C] = 8'h00;
mem[16'hA76D] = 8'hA7;
mem[16'hA76E] = 8'h00;
mem[16'hA76F] = 8'h9A;
mem[16'hA770] = 8'h00;
mem[16'hA771] = 8'hF0;
mem[16'hA772] = 8'h00;
mem[16'hA773] = 8'h20;
mem[16'hA774] = 8'h00;
mem[16'hA775] = 8'hA7;
mem[16'hA776] = 8'h00;
mem[16'hA777] = 8'h0A;
mem[16'hA778] = 8'h00;
mem[16'hA779] = 8'h40;
mem[16'hA77A] = 8'h00;
mem[16'hA77B] = 8'h44;
mem[16'hA77C] = 8'h00;
mem[16'hA77D] = 8'h41;
mem[16'hA77E] = 8'h00;
mem[16'hA77F] = 8'h45;
mem[16'hA780] = 8'h00;
mem[16'hA781] = 8'hEC;
mem[16'hA782] = 8'h00;
mem[16'hA783] = 8'h1D;
mem[16'hA784] = 8'h00;
mem[16'hA785] = 8'h40;
mem[16'hA786] = 8'h00;
mem[16'hA787] = 8'h75;
mem[16'hA788] = 8'h00;
mem[16'hA789] = 8'hD0;
mem[16'hA78A] = 8'h00;
mem[16'hA78B] = 8'h88;
mem[16'hA78C] = 8'h00;
mem[16'hA78D] = 8'hF6;
mem[16'hA78E] = 8'h00;
mem[16'hA78F] = 8'h60;
mem[16'hA790] = 8'h00;
mem[16'hA791] = 8'h60;
mem[16'hA792] = 8'h00;
mem[16'hA793] = 8'h00;
mem[16'hA794] = 8'h00;
mem[16'hA795] = 8'hAE;
mem[16'hA796] = 8'h00;
mem[16'hA797] = 8'h9D;
mem[16'hA798] = 8'h00;
mem[16'hA799] = 8'h0A;
mem[16'hA79A] = 8'h00;
mem[16'hA79B] = 8'h25;
mem[16'hA79C] = 8'h00;
mem[16'hA79D] = 8'h40;
mem[16'hA79E] = 8'h00;
mem[16'hA79F] = 8'h09;
mem[16'hA7A0] = 8'h00;
mem[16'hA7A1] = 8'h88;
mem[16'hA7A2] = 8'h00;
mem[16'hA7A3] = 8'h40;
mem[16'hA7A4] = 8'h00;
mem[16'hA7A5] = 8'h41;
mem[16'hA7A6] = 8'h00;
mem[16'hA7A7] = 8'h40;
mem[16'hA7A8] = 8'h00;
mem[16'hA7A9] = 8'h60;
mem[16'hA7AA] = 8'h00;
mem[16'hA7AB] = 8'h00;
mem[16'hA7AC] = 8'h00;
mem[16'hA7AD] = 8'h40;
mem[16'hA7AE] = 8'h00;
mem[16'hA7AF] = 8'hAD;
mem[16'hA7B0] = 8'h00;
mem[16'hA7B1] = 8'hAA;
mem[16'hA7B2] = 8'h00;
mem[16'hA7B3] = 8'h0E;
mem[16'hA7B4] = 8'h00;
mem[16'hA7B5] = 8'hB4;
mem[16'hA7B6] = 8'h00;
mem[16'hA7B7] = 8'hC5;
mem[16'hA7B8] = 8'h00;
mem[16'hA7B9] = 8'hD0;
mem[16'hA7BA] = 8'h00;
mem[16'hA7BB] = 8'hAD;
mem[16'hA7BC] = 8'h00;
mem[16'hA7BD] = 8'hAA;
mem[16'hA7BE] = 8'h00;
mem[16'hA7BF] = 8'h41;
mem[16'hA7C0] = 8'h00;
mem[16'hA7C1] = 8'h01;
mem[16'hA7C2] = 8'h00;
mem[16'hA7C3] = 8'h60;
mem[16'hA7C4] = 8'h00;
mem[16'hA7C5] = 8'hC2;
mem[16'hA7C6] = 8'h00;
mem[16'hA7C7] = 8'hF0;
mem[16'hA7C8] = 8'h00;
mem[16'hA7C9] = 8'h29;
mem[16'hA7CA] = 8'h00;
mem[16'hA7CB] = 8'hF0;
mem[16'hA7CC] = 8'h00;
mem[16'hA7CD] = 8'h20;
mem[16'hA7CE] = 8'h00;
mem[16'hA7CF] = 8'hA2;
mem[16'hA7D0] = 8'h00;
mem[16'hA7D1] = 8'hD0;
mem[16'hA7D2] = 8'h00;
mem[16'hA7D3] = 8'h60;
mem[16'hA7D4] = 8'h00;
mem[16'hA7D5] = 8'hAD;
mem[16'hA7D6] = 8'h00;
mem[16'hA7D7] = 8'h9D;
mem[16'hA7D8] = 8'h00;
mem[16'hA7D9] = 8'h40;
mem[16'hA7DA] = 8'h00;
mem[16'hA7DB] = 8'h01;
mem[16'hA7DC] = 8'h00;
mem[16'hA7DD] = 8'h85;
mem[16'hA7DE] = 8'h00;
mem[16'hA7DF] = 8'hAD;
mem[16'hA7E0] = 8'h00;
mem[16'hA7E1] = 8'hAA;
mem[16'hA7E2] = 8'h00;
mem[16'hA7E3] = 8'h63;
mem[16'hA7E4] = 8'h00;
mem[16'hA7E5] = 8'hA0;
mem[16'hA7E6] = 8'h00;
mem[16'hA7E7] = 8'h98;
mem[16'hA7E8] = 8'h00;
mem[16'hA7E9] = 8'h40;
mem[16'hA7EA] = 8'h00;
mem[16'hA7EB] = 8'h1E;
mem[16'hA7EC] = 8'h00;
mem[16'hA7ED] = 8'hA5;
mem[16'hA7EE] = 8'h00;
mem[16'hA7EF] = 8'hE9;
mem[16'hA7F0] = 8'h00;
mem[16'hA7F1] = 8'h91;
mem[16'hA7F2] = 8'h00;
mem[16'hA7F3] = 8'h48;
mem[16'hA7F4] = 8'h00;
mem[16'hA7F5] = 8'h41;
mem[16'hA7F6] = 8'h00;
mem[16'hA7F7] = 8'h00;
mem[16'hA7F8] = 8'h00;
mem[16'hA7F9] = 8'h91;
mem[16'hA7FA] = 8'h00;
mem[16'hA7FB] = 8'hAA;
mem[16'hA7FC] = 8'h00;
mem[16'hA7FD] = 8'h68;
mem[16'hA7FE] = 8'h00;
mem[16'hA7FF] = 8'hC8;
mem[16'hA800] = 8'h85;
mem[16'hA801] = 8'hA9;
mem[16'hA802] = 8'hB3;
mem[16'hA803] = 8'h48;
mem[16'hA804] = 8'hA9;
mem[16'hA805] = 8'hFF;
mem[16'hA806] = 8'h48;
mem[16'hA807] = 8'h60;
mem[16'hA808] = 8'h02;
mem[16'hA809] = 8'h02;
mem[16'hA80A] = 8'h02;
mem[16'hA80B] = 8'h02;
mem[16'hA80C] = 8'h02;
mem[16'hA80D] = 8'h02;
mem[16'hA80E] = 8'h02;
mem[16'hA80F] = 8'h02;
mem[16'hA810] = 8'h02;
mem[16'hA811] = 8'h02;
mem[16'hA812] = 8'h02;
mem[16'hA813] = 8'h02;
mem[16'hA814] = 8'h02;
mem[16'hA815] = 8'h02;
mem[16'hA816] = 8'h02;
mem[16'hA817] = 8'h02;
mem[16'hA818] = 8'h02;
mem[16'hA819] = 8'h02;
mem[16'hA81A] = 8'h02;
mem[16'hA81B] = 8'h02;
mem[16'hA81C] = 8'h02;
mem[16'hA81D] = 8'h02;
mem[16'hA81E] = 8'h02;
mem[16'hA81F] = 8'h02;
mem[16'hA820] = 8'h02;
mem[16'hA821] = 8'h02;
mem[16'hA822] = 8'h02;
mem[16'hA823] = 8'h02;
mem[16'hA824] = 8'h81;
mem[16'hA825] = 8'h81;
mem[16'hA826] = 8'h81;
mem[16'hA827] = 8'h81;
mem[16'hA828] = 8'h81;
mem[16'hA829] = 8'h81;
mem[16'hA82A] = 8'h81;
mem[16'hA82B] = 8'h81;
mem[16'hA82C] = 8'h81;
mem[16'hA82D] = 8'h81;
mem[16'hA82E] = 8'h81;
mem[16'hA82F] = 8'h81;
mem[16'hA830] = 8'h81;
mem[16'hA831] = 8'h81;
mem[16'hA832] = 8'h81;
mem[16'hA833] = 8'h81;
mem[16'hA834] = 8'h81;
mem[16'hA835] = 8'h81;
mem[16'hA836] = 8'h81;
mem[16'hA837] = 8'h81;
mem[16'hA838] = 8'h81;
mem[16'hA839] = 8'h81;
mem[16'hA83A] = 8'h81;
mem[16'hA83B] = 8'h81;
mem[16'hA83C] = 8'h81;
mem[16'hA83D] = 8'h81;
mem[16'hA83E] = 8'h81;
mem[16'hA83F] = 8'h81;
mem[16'hA840] = 8'h81;
mem[16'hA841] = 8'h81;
mem[16'hA842] = 8'h81;
mem[16'hA843] = 8'h81;
mem[16'hA844] = 8'h81;
mem[16'hA845] = 8'h81;
mem[16'hA846] = 8'h81;
mem[16'hA847] = 8'h81;
mem[16'hA848] = 8'h81;
mem[16'hA849] = 8'h81;
mem[16'hA84A] = 8'h81;
mem[16'hA84B] = 8'h81;
mem[16'hA84C] = 8'h81;
mem[16'hA84D] = 8'h81;
mem[16'hA84E] = 8'h81;
mem[16'hA84F] = 8'h81;
mem[16'hA850] = 8'h81;
mem[16'hA851] = 8'h81;
mem[16'hA852] = 8'h81;
mem[16'hA853] = 8'h81;
mem[16'hA854] = 8'h81;
mem[16'hA855] = 8'h81;
mem[16'hA856] = 8'h81;
mem[16'hA857] = 8'h81;
mem[16'hA858] = 8'h81;
mem[16'hA859] = 8'h81;
mem[16'hA85A] = 8'h81;
mem[16'hA85B] = 8'h81;
mem[16'hA85C] = 8'h81;
mem[16'hA85D] = 8'h81;
mem[16'hA85E] = 8'h81;
mem[16'hA85F] = 8'h81;
mem[16'hA860] = 8'h81;
mem[16'hA861] = 8'h81;
mem[16'hA862] = 8'h81;
mem[16'hA863] = 8'h81;
mem[16'hA864] = 8'h81;
mem[16'hA865] = 8'h81;
mem[16'hA866] = 8'h81;
mem[16'hA867] = 8'h81;
mem[16'hA868] = 8'h81;
mem[16'hA869] = 8'h81;
mem[16'hA86A] = 8'h81;
mem[16'hA86B] = 8'h81;
mem[16'hA86C] = 8'h81;
mem[16'hA86D] = 8'h81;
mem[16'hA86E] = 8'h81;
mem[16'hA86F] = 8'h81;
mem[16'hA870] = 8'h81;
mem[16'hA871] = 8'h81;
mem[16'hA872] = 8'h81;
mem[16'hA873] = 8'h81;
mem[16'hA874] = 8'h81;
mem[16'hA875] = 8'h81;
mem[16'hA876] = 8'h81;
mem[16'hA877] = 8'h81;
mem[16'hA878] = 8'h81;
mem[16'hA879] = 8'h81;
mem[16'hA87A] = 8'h81;
mem[16'hA87B] = 8'h81;
mem[16'hA87C] = 8'h81;
mem[16'hA87D] = 8'h81;
mem[16'hA87E] = 8'h81;
mem[16'hA87F] = 8'h81;
mem[16'hA880] = 8'h81;
mem[16'hA881] = 8'h81;
mem[16'hA882] = 8'h81;
mem[16'hA883] = 8'h81;
mem[16'hA884] = 8'h81;
mem[16'hA885] = 8'h81;
mem[16'hA886] = 8'h81;
mem[16'hA887] = 8'h81;
mem[16'hA888] = 8'h81;
mem[16'hA889] = 8'h81;
mem[16'hA88A] = 8'h81;
mem[16'hA88B] = 8'h81;
mem[16'hA88C] = 8'h53;
mem[16'hA88D] = 8'h41;
mem[16'hA88E] = 8'h56;
mem[16'hA88F] = 8'hC5;
mem[16'hA890] = 8'h52;
mem[16'hA891] = 8'h55;
mem[16'hA892] = 8'hCE;
mem[16'hA893] = 8'h43;
mem[16'hA894] = 8'h48;
mem[16'hA895] = 8'h41;
mem[16'hA896] = 8'h49;
mem[16'hA897] = 8'hCE;
mem[16'hA898] = 8'h44;
mem[16'hA899] = 8'h45;
mem[16'hA89A] = 8'h4C;
mem[16'hA89B] = 8'h45;
mem[16'hA89C] = 8'h54;
mem[16'hA89D] = 8'hC5;
mem[16'hA89E] = 8'h4C;
mem[16'hA89F] = 8'h4F;
mem[16'hA8A0] = 8'h43;
mem[16'hA8A1] = 8'hCB;
mem[16'hA8A2] = 8'h55;
mem[16'hA8A3] = 8'h4E;
mem[16'hA8A4] = 8'h4C;
mem[16'hA8A5] = 8'h4F;
mem[16'hA8A6] = 8'h43;
mem[16'hA8A7] = 8'hCB;
mem[16'hA8A8] = 8'h43;
mem[16'hA8A9] = 8'h4C;
mem[16'hA8AA] = 8'h4F;
mem[16'hA8AB] = 8'h53;
mem[16'hA8AC] = 8'hC5;
mem[16'hA8AD] = 8'h52;
mem[16'hA8AE] = 8'h45;
mem[16'hA8AF] = 8'h41;
mem[16'hA8B0] = 8'hC4;
mem[16'hA8B1] = 8'h45;
mem[16'hA8B2] = 8'h58;
mem[16'hA8B3] = 8'h45;
mem[16'hA8B4] = 8'hC3;
mem[16'hA8B5] = 8'h57;
mem[16'hA8B6] = 8'h52;
mem[16'hA8B7] = 8'h49;
mem[16'hA8B8] = 8'h54;
mem[16'hA8B9] = 8'hC5;
mem[16'hA8BA] = 8'h50;
mem[16'hA8BB] = 8'h4F;
mem[16'hA8BC] = 8'h53;
mem[16'hA8BD] = 8'h49;
mem[16'hA8BE] = 8'h54;
mem[16'hA8BF] = 8'h49;
mem[16'hA8C0] = 8'h4F;
mem[16'hA8C1] = 8'hCE;
mem[16'hA8C2] = 8'h4F;
mem[16'hA8C3] = 8'h50;
mem[16'hA8C4] = 8'h45;
mem[16'hA8C5] = 8'hCE;
mem[16'hA8C6] = 8'h41;
mem[16'hA8C7] = 8'h50;
mem[16'hA8C8] = 8'h50;
mem[16'hA8C9] = 8'h45;
mem[16'hA8CA] = 8'h4E;
mem[16'hA8CB] = 8'hC4;
mem[16'hA8CC] = 8'h52;
mem[16'hA8CD] = 8'h45;
mem[16'hA8CE] = 8'h4E;
mem[16'hA8CF] = 8'h41;
mem[16'hA8D0] = 8'h4D;
mem[16'hA8D1] = 8'hC5;
mem[16'hA8D2] = 8'h43;
mem[16'hA8D3] = 8'h41;
mem[16'hA8D4] = 8'h54;
mem[16'hA8D5] = 8'h41;
mem[16'hA8D6] = 8'h4C;
mem[16'hA8D7] = 8'h4F;
mem[16'hA8D8] = 8'hC7;
mem[16'hA8D9] = 8'h4D;
mem[16'hA8DA] = 8'h4F;
mem[16'hA8DB] = 8'hCE;
mem[16'hA8DC] = 8'h4E;
mem[16'hA8DD] = 8'h4F;
mem[16'hA8DE] = 8'h4D;
mem[16'hA8DF] = 8'h4F;
mem[16'hA8E0] = 8'hCE;
mem[16'hA8E1] = 8'h50;
mem[16'hA8E2] = 8'h52;
mem[16'hA8E3] = 8'hA3;
mem[16'hA8E4] = 8'h49;
mem[16'hA8E5] = 8'h4E;
mem[16'hA8E6] = 8'hA3;
mem[16'hA8E7] = 8'h4D;
mem[16'hA8E8] = 8'h41;
mem[16'hA8E9] = 8'h58;
mem[16'hA8EA] = 8'h46;
mem[16'hA8EB] = 8'h49;
mem[16'hA8EC] = 8'h4C;
mem[16'hA8ED] = 8'h45;
mem[16'hA8EE] = 8'hD3;
mem[16'hA8EF] = 8'h46;
mem[16'hA8F0] = 8'hD0;
mem[16'hA8F1] = 8'h49;
mem[16'hA8F2] = 8'h4E;
mem[16'hA8F3] = 8'hD4;
mem[16'hA8F4] = 8'h42;
mem[16'hA8F5] = 8'h53;
mem[16'hA8F6] = 8'h41;
mem[16'hA8F7] = 8'h56;
mem[16'hA8F8] = 8'hC5;
mem[16'hA8F9] = 8'h42;
mem[16'hA8FA] = 8'h4C;
mem[16'hA8FB] = 8'h4F;
mem[16'hA8FC] = 8'h41;
mem[16'hA8FD] = 8'hC4;
mem[16'hA8FE] = 8'h42;
mem[16'hA8FF] = 8'h52;
mem[16'hA900] = 8'h20;
mem[16'hA901] = 8'h21;
mem[16'hA902] = 8'h22;
mem[16'hA903] = 8'h23;
mem[16'hA904] = 8'h24;
mem[16'hA905] = 8'h25;
mem[16'hA906] = 8'h26;
mem[16'hA907] = 8'h27;
mem[16'hA908] = 8'h28;
mem[16'hA909] = 8'h29;
mem[16'hA90A] = 8'h2A;
mem[16'hA90B] = 8'h2B;
mem[16'hA90C] = 8'h2C;
mem[16'hA90D] = 8'h2D;
mem[16'hA90E] = 8'h2E;
mem[16'hA90F] = 8'h2F;
mem[16'hA910] = 8'h30;
mem[16'hA911] = 8'h31;
mem[16'hA912] = 8'h32;
mem[16'hA913] = 8'h33;
mem[16'hA914] = 8'h34;
mem[16'hA915] = 8'h35;
mem[16'hA916] = 8'h36;
mem[16'hA917] = 8'h37;
mem[16'hA918] = 8'h38;
mem[16'hA919] = 8'h39;
mem[16'hA91A] = 8'h3A;
mem[16'hA91B] = 8'h3B;
mem[16'hA91C] = 8'h3C;
mem[16'hA91D] = 8'h3D;
mem[16'hA91E] = 8'h3E;
mem[16'hA91F] = 8'h3F;
mem[16'hA920] = 8'hFF;
mem[16'hA921] = 8'h61;
mem[16'hA922] = 8'h62;
mem[16'hA923] = 8'h63;
mem[16'hA924] = 8'h64;
mem[16'hA925] = 8'h65;
mem[16'hA926] = 8'h66;
mem[16'hA927] = 8'h67;
mem[16'hA928] = 8'h68;
mem[16'hA929] = 8'h69;
mem[16'hA92A] = 8'h6A;
mem[16'hA92B] = 8'h6B;
mem[16'hA92C] = 8'h6C;
mem[16'hA92D] = 8'h6D;
mem[16'hA92E] = 8'h6E;
mem[16'hA92F] = 8'h6F;
mem[16'hA930] = 8'h70;
mem[16'hA931] = 8'h71;
mem[16'hA932] = 8'h72;
mem[16'hA933] = 8'h73;
mem[16'hA934] = 8'h74;
mem[16'hA935] = 8'h75;
mem[16'hA936] = 8'h76;
mem[16'hA937] = 8'h77;
mem[16'hA938] = 8'h78;
mem[16'hA939] = 8'h79;
mem[16'hA93A] = 8'h7A;
mem[16'hA93B] = 8'h7B;
mem[16'hA93C] = 8'h7C;
mem[16'hA93D] = 8'h7D;
mem[16'hA93E] = 8'h7E;
mem[16'hA93F] = 8'h7F;
mem[16'hA940] = 8'h80;
mem[16'hA941] = 8'h81;
mem[16'hA942] = 8'h82;
mem[16'hA943] = 8'h83;
mem[16'hA944] = 8'h84;
mem[16'hA945] = 8'h85;
mem[16'hA946] = 8'h86;
mem[16'hA947] = 8'h87;
mem[16'hA948] = 8'h88;
mem[16'hA949] = 8'h89;
mem[16'hA94A] = 8'h8A;
mem[16'hA94B] = 8'h8B;
mem[16'hA94C] = 8'h8C;
mem[16'hA94D] = 8'h8D;
mem[16'hA94E] = 8'h8E;
mem[16'hA94F] = 8'h8F;
mem[16'hA950] = 8'h90;
mem[16'hA951] = 8'h91;
mem[16'hA952] = 8'h92;
mem[16'hA953] = 8'h93;
mem[16'hA954] = 8'h94;
mem[16'hA955] = 8'h95;
mem[16'hA956] = 8'h96;
mem[16'hA957] = 8'h97;
mem[16'hA958] = 8'h98;
mem[16'hA959] = 8'h99;
mem[16'hA95A] = 8'h9A;
mem[16'hA95B] = 8'h9B;
mem[16'hA95C] = 8'h9C;
mem[16'hA95D] = 8'h9D;
mem[16'hA95E] = 8'h9E;
mem[16'hA95F] = 8'h9F;
mem[16'hA960] = 8'hFF;
mem[16'hA961] = 8'h01;
mem[16'hA962] = 8'h00;
mem[16'hA963] = 8'hFF;
mem[16'hA964] = 8'h7F;
mem[16'hA965] = 8'h00;
mem[16'hA966] = 8'h00;
mem[16'hA967] = 8'hFF;
mem[16'hA968] = 8'h7F;
mem[16'hA969] = 8'h00;
mem[16'hA96A] = 8'h00;
mem[16'hA96B] = 8'hFF;
mem[16'hA96C] = 8'h7F;
mem[16'hA96D] = 8'h00;
mem[16'hA96E] = 8'h00;
mem[16'hA96F] = 8'hFF;
mem[16'hA970] = 8'hFF;
mem[16'hA971] = 8'h0D;
mem[16'hA972] = 8'h07;
mem[16'hA973] = 8'h8D;
mem[16'hA974] = 8'h4C;
mem[16'hA975] = 8'h41;
mem[16'hA976] = 8'h4E;
mem[16'hA977] = 8'h47;
mem[16'hA978] = 8'h55;
mem[16'hA979] = 8'h41;
mem[16'hA97A] = 8'h47;
mem[16'hA97B] = 8'h45;
mem[16'hA97C] = 8'h20;
mem[16'hA97D] = 8'h4E;
mem[16'hA97E] = 8'h4F;
mem[16'hA97F] = 8'h54;
mem[16'hA980] = 8'h20;
mem[16'hA981] = 8'h41;
mem[16'hA982] = 8'h56;
mem[16'hA983] = 8'h41;
mem[16'hA984] = 8'h49;
mem[16'hA985] = 8'h4C;
mem[16'hA986] = 8'h41;
mem[16'hA987] = 8'h42;
mem[16'hA988] = 8'h4C;
mem[16'hA989] = 8'hC5;
mem[16'hA98A] = 8'h52;
mem[16'hA98B] = 8'h41;
mem[16'hA98C] = 8'h4E;
mem[16'hA98D] = 8'h47;
mem[16'hA98E] = 8'h45;
mem[16'hA98F] = 8'h20;
mem[16'hA990] = 8'h45;
mem[16'hA991] = 8'h52;
mem[16'hA992] = 8'h52;
mem[16'hA993] = 8'h4F;
mem[16'hA994] = 8'hD2;
mem[16'hA995] = 8'h57;
mem[16'hA996] = 8'h52;
mem[16'hA997] = 8'h49;
mem[16'hA998] = 8'h54;
mem[16'hA999] = 8'h45;
mem[16'hA99A] = 8'h20;
mem[16'hA99B] = 8'h50;
mem[16'hA99C] = 8'h52;
mem[16'hA99D] = 8'h4F;
mem[16'hA99E] = 8'h54;
mem[16'hA99F] = 8'h45;
mem[16'hA9A0] = 8'h43;
mem[16'hA9A1] = 8'h54;
mem[16'hA9A2] = 8'h45;
mem[16'hA9A3] = 8'hC4;
mem[16'hA9A4] = 8'h45;
mem[16'hA9A5] = 8'h4E;
mem[16'hA9A6] = 8'h44;
mem[16'hA9A7] = 8'h20;
mem[16'hA9A8] = 8'h4F;
mem[16'hA9A9] = 8'h46;
mem[16'hA9AA] = 8'h20;
mem[16'hA9AB] = 8'h44;
mem[16'hA9AC] = 8'h41;
mem[16'hA9AD] = 8'h54;
mem[16'hA9AE] = 8'hC1;
mem[16'hA9AF] = 8'h46;
mem[16'hA9B0] = 8'h49;
mem[16'hA9B1] = 8'h4C;
mem[16'hA9B2] = 8'h45;
mem[16'hA9B3] = 8'h20;
mem[16'hA9B4] = 8'h4E;
mem[16'hA9B5] = 8'h4F;
mem[16'hA9B6] = 8'h54;
mem[16'hA9B7] = 8'h20;
mem[16'hA9B8] = 8'h46;
mem[16'hA9B9] = 8'h4F;
mem[16'hA9BA] = 8'h55;
mem[16'hA9BB] = 8'h4E;
mem[16'hA9BC] = 8'hC4;
mem[16'hA9BD] = 8'h56;
mem[16'hA9BE] = 8'h4F;
mem[16'hA9BF] = 8'h4C;
mem[16'hA9C0] = 8'h55;
mem[16'hA9C1] = 8'h4D;
mem[16'hA9C2] = 8'h45;
mem[16'hA9C3] = 8'h20;
mem[16'hA9C4] = 8'h4D;
mem[16'hA9C5] = 8'h49;
mem[16'hA9C6] = 8'h53;
mem[16'hA9C7] = 8'h4D;
mem[16'hA9C8] = 8'h41;
mem[16'hA9C9] = 8'h54;
mem[16'hA9CA] = 8'h43;
mem[16'hA9CB] = 8'hC8;
mem[16'hA9CC] = 8'h49;
mem[16'hA9CD] = 8'h2F;
mem[16'hA9CE] = 8'h4F;
mem[16'hA9CF] = 8'h20;
mem[16'hA9D0] = 8'h45;
mem[16'hA9D1] = 8'h52;
mem[16'hA9D2] = 8'h52;
mem[16'hA9D3] = 8'h4F;
mem[16'hA9D4] = 8'hD2;
mem[16'hA9D5] = 8'h44;
mem[16'hA9D6] = 8'h49;
mem[16'hA9D7] = 8'h53;
mem[16'hA9D8] = 8'h4B;
mem[16'hA9D9] = 8'h20;
mem[16'hA9DA] = 8'h46;
mem[16'hA9DB] = 8'h55;
mem[16'hA9DC] = 8'h4C;
mem[16'hA9DD] = 8'hCC;
mem[16'hA9DE] = 8'h46;
mem[16'hA9DF] = 8'h49;
mem[16'hA9E0] = 8'h4C;
mem[16'hA9E1] = 8'h45;
mem[16'hA9E2] = 8'h20;
mem[16'hA9E3] = 8'h4C;
mem[16'hA9E4] = 8'h4F;
mem[16'hA9E5] = 8'h43;
mem[16'hA9E6] = 8'h4B;
mem[16'hA9E7] = 8'h45;
mem[16'hA9E8] = 8'hC4;
mem[16'hA9E9] = 8'h53;
mem[16'hA9EA] = 8'h59;
mem[16'hA9EB] = 8'h4E;
mem[16'hA9EC] = 8'h54;
mem[16'hA9ED] = 8'h41;
mem[16'hA9EE] = 8'h58;
mem[16'hA9EF] = 8'h20;
mem[16'hA9F0] = 8'h45;
mem[16'hA9F1] = 8'h52;
mem[16'hA9F2] = 8'h52;
mem[16'hA9F3] = 8'h4F;
mem[16'hA9F4] = 8'hD2;
mem[16'hA9F5] = 8'h4E;
mem[16'hA9F6] = 8'h4F;
mem[16'hA9F7] = 8'h20;
mem[16'hA9F8] = 8'h42;
mem[16'hA9F9] = 8'h55;
mem[16'hA9FA] = 8'h46;
mem[16'hA9FB] = 8'h46;
mem[16'hA9FC] = 8'h45;
mem[16'hA9FD] = 8'h52;
mem[16'hA9FE] = 8'h53;
mem[16'hA9FF] = 8'h20;
mem[16'hAA00] = 8'h04;
mem[16'hAA01] = 8'h04;
mem[16'hAA02] = 8'h04;
mem[16'hAA03] = 8'h04;
mem[16'hAA04] = 8'h05;
mem[16'hAA05] = 8'h05;
mem[16'hAA06] = 8'h05;
mem[16'hAA07] = 8'h05;
mem[16'hAA08] = 8'h06;
mem[16'hAA09] = 8'h06;
mem[16'hAA0A] = 8'h06;
mem[16'hAA0B] = 8'h06;
mem[16'hAA0C] = 8'h07;
mem[16'hAA0D] = 8'h07;
mem[16'hAA0E] = 8'h07;
mem[16'hAA0F] = 8'h07;
mem[16'hAA10] = 8'h08;
mem[16'hAA11] = 8'h08;
mem[16'hAA12] = 8'h08;
mem[16'hAA13] = 8'h08;
mem[16'hAA14] = 8'h09;
mem[16'hAA15] = 8'h09;
mem[16'hAA16] = 8'h09;
mem[16'hAA17] = 8'h09;
mem[16'hAA18] = 8'h0A;
mem[16'hAA19] = 8'h0A;
mem[16'hAA1A] = 8'h0A;
mem[16'hAA1B] = 8'h0A;
mem[16'hAA1C] = 8'h0B;
mem[16'hAA1D] = 8'h0B;
mem[16'hAA1E] = 8'h0B;
mem[16'hAA1F] = 8'h0B;
mem[16'hAA20] = 8'hFF;
mem[16'hAA21] = 8'h14;
mem[16'hAA22] = 8'h14;
mem[16'hAA23] = 8'h14;
mem[16'hAA24] = 8'h15;
mem[16'hAA25] = 8'h15;
mem[16'hAA26] = 8'h15;
mem[16'hAA27] = 8'h15;
mem[16'hAA28] = 8'h16;
mem[16'hAA29] = 8'h16;
mem[16'hAA2A] = 8'h16;
mem[16'hAA2B] = 8'h16;
mem[16'hAA2C] = 8'h17;
mem[16'hAA2D] = 8'h17;
mem[16'hAA2E] = 8'h17;
mem[16'hAA2F] = 8'h17;
mem[16'hAA30] = 8'h18;
mem[16'hAA31] = 8'h18;
mem[16'hAA32] = 8'h18;
mem[16'hAA33] = 8'h18;
mem[16'hAA34] = 8'h19;
mem[16'hAA35] = 8'h19;
mem[16'hAA36] = 8'h19;
mem[16'hAA37] = 8'h19;
mem[16'hAA38] = 8'h1A;
mem[16'hAA39] = 8'h1A;
mem[16'hAA3A] = 8'h1A;
mem[16'hAA3B] = 8'h1A;
mem[16'hAA3C] = 8'h1B;
mem[16'hAA3D] = 8'h1B;
mem[16'hAA3E] = 8'h1B;
mem[16'hAA3F] = 8'h1B;
mem[16'hAA40] = 8'h1C;
mem[16'hAA41] = 8'h1C;
mem[16'hAA42] = 8'h1C;
mem[16'hAA43] = 8'h1C;
mem[16'hAA44] = 8'h1D;
mem[16'hAA45] = 8'h1D;
mem[16'hAA46] = 8'h1D;
mem[16'hAA47] = 8'h1D;
mem[16'hAA48] = 8'h1E;
mem[16'hAA49] = 8'h1E;
mem[16'hAA4A] = 8'h1E;
mem[16'hAA4B] = 8'h1E;
mem[16'hAA4C] = 8'h1F;
mem[16'hAA4D] = 8'h1F;
mem[16'hAA4E] = 8'h1F;
mem[16'hAA4F] = 8'h1F;
mem[16'hAA50] = 8'h20;
mem[16'hAA51] = 8'h20;
mem[16'hAA52] = 8'h20;
mem[16'hAA53] = 8'h20;
mem[16'hAA54] = 8'h21;
mem[16'hAA55] = 8'h21;
mem[16'hAA56] = 8'h21;
mem[16'hAA57] = 8'h21;
mem[16'hAA58] = 8'h22;
mem[16'hAA59] = 8'h22;
mem[16'hAA5A] = 8'h22;
mem[16'hAA5B] = 8'h22;
mem[16'hAA5C] = 8'h23;
mem[16'hAA5D] = 8'h23;
mem[16'hAA5E] = 8'h23;
mem[16'hAA5F] = 8'h23;
mem[16'hAA60] = 8'hFF;
mem[16'hAA61] = 8'h00;
mem[16'hAA62] = 8'h00;
mem[16'hAA63] = 8'h06;
mem[16'hAA64] = 8'h03;
mem[16'hAA65] = 8'h00;
mem[16'hAA66] = 8'hFE;
mem[16'hAA67] = 8'h00;
mem[16'hAA68] = 8'h01;
mem[16'hAA69] = 8'h00;
mem[16'hAA6A] = 8'h06;
mem[16'hAA6B] = 8'h00;
mem[16'hAA6C] = 8'h01;
mem[16'hAA6D] = 8'h00;
mem[16'hAA6E] = 8'h00;
mem[16'hAA6F] = 8'h00;
mem[16'hAA70] = 8'h00;
mem[16'hAA71] = 8'h00;
mem[16'hAA72] = 8'h00;
mem[16'hAA73] = 8'h40;
mem[16'hAA74] = 8'h00;
mem[16'hAA75] = 8'h00;
mem[16'hAA76] = 8'hAE;
mem[16'hAA77] = 8'hA4;
mem[16'hAA78] = 8'hB4;
mem[16'hAA79] = 8'hB0;
mem[16'hAA7A] = 8'hAD;
mem[16'hAA7B] = 8'hA4;
mem[16'hAA7C] = 8'hB9;
mem[16'hAA7D] = 8'hB6;
mem[16'hAA7E] = 8'hA0;
mem[16'hAA7F] = 8'hA0;
mem[16'hAA80] = 8'hA0;
mem[16'hAA81] = 8'hA0;
mem[16'hAA82] = 8'hA0;
mem[16'hAA83] = 8'hA0;
mem[16'hAA84] = 8'hA0;
mem[16'hAA85] = 8'hA0;
mem[16'hAA86] = 8'hA0;
mem[16'hAA87] = 8'hA0;
mem[16'hAA88] = 8'hA0;
mem[16'hAA89] = 8'hA0;
mem[16'hAA8A] = 8'hA0;
mem[16'hAA8B] = 8'hA0;
mem[16'hAA8C] = 8'hA0;
mem[16'hAA8D] = 8'hA0;
mem[16'hAA8E] = 8'hA0;
mem[16'hAA8F] = 8'hA0;
mem[16'hAA90] = 8'hA0;
mem[16'hAA91] = 8'hA0;
mem[16'hAA92] = 8'hA0;
mem[16'hAA93] = 8'hA0;
mem[16'hAA94] = 8'hA0;
mem[16'hAA95] = 8'hA0;
mem[16'hAA96] = 8'hA0;
mem[16'hAA97] = 8'hA0;
mem[16'hAA98] = 8'hA0;
mem[16'hAA99] = 8'hA0;
mem[16'hAA9A] = 8'hA0;
mem[16'hAA9B] = 8'hA0;
mem[16'hAA9C] = 8'hA0;
mem[16'hAA9D] = 8'hA0;
mem[16'hAA9E] = 8'hA0;
mem[16'hAA9F] = 8'hA0;
mem[16'hAAA0] = 8'hA0;
mem[16'hAAA1] = 8'hA0;
mem[16'hAAA2] = 8'hA0;
mem[16'hAAA3] = 8'hA0;
mem[16'hAAA4] = 8'hA0;
mem[16'hAAA5] = 8'hA0;
mem[16'hAAA6] = 8'hA0;
mem[16'hAAA7] = 8'hA0;
mem[16'hAAA8] = 8'hA0;
mem[16'hAAA9] = 8'hA0;
mem[16'hAAAA] = 8'hA0;
mem[16'hAAAB] = 8'hA0;
mem[16'hAAAC] = 8'hA0;
mem[16'hAAAD] = 8'hA0;
mem[16'hAAAE] = 8'hA0;
mem[16'hAAAF] = 8'hA0;
mem[16'hAAB0] = 8'hA0;
mem[16'hAAB1] = 8'h03;
mem[16'hAAB2] = 8'h84;
mem[16'hAAB3] = 8'h00;
mem[16'hAAB4] = 8'h00;
mem[16'hAAB5] = 8'h00;
mem[16'hAAB6] = 8'h40;
mem[16'hAAB7] = 8'h00;
mem[16'hAAB8] = 8'hC1;
mem[16'hAAB9] = 8'hD0;
mem[16'hAABA] = 8'hD0;
mem[16'hAABB] = 8'hCC;
mem[16'hAABC] = 8'hC5;
mem[16'hAABD] = 8'hD3;
mem[16'hAABE] = 8'hCF;
mem[16'hAABF] = 8'hC6;
mem[16'hAAC0] = 8'hD4;
mem[16'hAAC1] = 8'hE8;
mem[16'hAAC2] = 8'hB7;
mem[16'hAAC3] = 8'hBB;
mem[16'hAAC4] = 8'hB3;
mem[16'hAAC5] = 8'hBB;
mem[16'hAAC6] = 8'hB4;
mem[16'hAAC7] = 8'h00;
mem[16'hAAC8] = 8'hC0;
mem[16'hAAC9] = 8'h7E;
mem[16'hAACA] = 8'hB3;
mem[16'hAACB] = 8'h21;
mem[16'hAACC] = 8'hAB;
mem[16'hAACD] = 8'h05;
mem[16'hAACE] = 8'hAC;
mem[16'hAACF] = 8'h57;
mem[16'hAAD0] = 8'hAC;
mem[16'hAAD1] = 8'h6F;
mem[16'hAAD2] = 8'hAC;
mem[16'hAAD3] = 8'h2A;
mem[16'hAAD4] = 8'hAD;
mem[16'hAAD5] = 8'h97;
mem[16'hAAD6] = 8'hAD;
mem[16'hAAD7] = 8'hEE;
mem[16'hAAD8] = 8'hAC;
mem[16'hAAD9] = 8'hF5;
mem[16'hAADA] = 8'hAC;
mem[16'hAADB] = 8'h39;
mem[16'hAADC] = 8'hAC;
mem[16'hAADD] = 8'h11;
mem[16'hAADE] = 8'hAD;
mem[16'hAADF] = 8'h8D;
mem[16'hAAE0] = 8'hAE;
mem[16'hAAE1] = 8'h17;
mem[16'hAAE2] = 8'hAD;
mem[16'hAAE3] = 8'h7E;
mem[16'hAAE4] = 8'hB3;
mem[16'hAAE5] = 8'h7E;
mem[16'hAAE6] = 8'hB3;
mem[16'hAAE7] = 8'h89;
mem[16'hAAE8] = 8'hAC;
mem[16'hAAE9] = 8'h95;
mem[16'hAAEA] = 8'hAC;
mem[16'hAAEB] = 8'h86;
mem[16'hAAEC] = 8'hAC;
mem[16'hAAED] = 8'h92;
mem[16'hAAEE] = 8'hAC;
mem[16'hAAEF] = 8'h7E;
mem[16'hAAF0] = 8'hB3;
mem[16'hAAF1] = 8'h7E;
mem[16'hAAF2] = 8'hB3;
mem[16'hAAF3] = 8'hBD;
mem[16'hAAF4] = 8'hAC;
mem[16'hAAF5] = 8'hC9;
mem[16'hAAF6] = 8'hAC;
mem[16'hAAF7] = 8'hBA;
mem[16'hAAF8] = 8'hAC;
mem[16'hAAF9] = 8'hC6;
mem[16'hAAFA] = 8'hAC;
mem[16'hAAFB] = 8'h7E;
mem[16'hAAFC] = 8'hB3;
mem[16'hAAFD] = 8'hE0;
mem[16'hAAFE] = 8'h00;
mem[16'hAAFF] = 8'hF0;
mem[16'hAB00] = 8'hAD;
mem[16'hAB01] = 8'hA9;
mem[16'hAB02] = 8'hB7;
mem[16'hAB03] = 8'hB3;
mem[16'hAB04] = 8'hAE;
mem[16'hAB05] = 8'hAA;
mem[16'hAB06] = 8'hB9;
mem[16'hAB07] = 8'hB4;
mem[16'hAB08] = 8'hAF;
mem[16'hAB09] = 8'hAB;
mem[16'hAB0A] = 8'hBA;
mem[16'hAB0B] = 8'hB5;
mem[16'hAB0C] = 8'hB2;
mem[16'hAB0D] = 8'hAC;
mem[16'hAB0E] = 8'hBB;
mem[16'hAB0F] = 8'hB6;
mem[16'hAB10] = 8'hB3;
mem[16'hAB11] = 8'hB7;
mem[16'hAB12] = 8'hA9;
mem[16'hAB13] = 8'hAD;
mem[16'hAB14] = 8'hB4;
mem[16'hAB15] = 8'hB9;
mem[16'hAB16] = 8'hAA;
mem[16'hAB17] = 8'hAE;
mem[16'hAB18] = 8'hB5;
mem[16'hAB19] = 8'hBA;
mem[16'hAB1A] = 8'hAB;
mem[16'hAB1B] = 8'hAF;
mem[16'hAB1C] = 8'hB6;
mem[16'hAB1D] = 8'hBB;
mem[16'hAB1E] = 8'hAC;
mem[16'hAB1F] = 8'hB2;
mem[16'hAB20] = 8'hFF;
mem[16'hAB21] = 8'hBC;
mem[16'hAB22] = 8'hD3;
mem[16'hAB23] = 8'hCD;
mem[16'hAB24] = 8'hCA;
mem[16'hAB25] = 8'hBD;
mem[16'hAB26] = 8'hD4;
mem[16'hAB27] = 8'hCE;
mem[16'hAB28] = 8'hCB;
mem[16'hAB29] = 8'hBE;
mem[16'hAB2A] = 8'hD5;
mem[16'hAB2B] = 8'hCF;
mem[16'hAB2C] = 8'hCC;
mem[16'hAB2D] = 8'hBF;
mem[16'hAB2E] = 8'hD6;
mem[16'hAB2F] = 8'hD2;
mem[16'hAB30] = 8'hCD;
mem[16'hAB31] = 8'hD3;
mem[16'hAB32] = 8'hBC;
mem[16'hAB33] = 8'hC9;
mem[16'hAB34] = 8'hCE;
mem[16'hAB35] = 8'hD4;
mem[16'hAB36] = 8'hBD;
mem[16'hAB37] = 8'hCA;
mem[16'hAB38] = 8'hCF;
mem[16'hAB39] = 8'hD5;
mem[16'hAB3A] = 8'hBE;
mem[16'hAB3B] = 8'hCB;
mem[16'hAB3C] = 8'hD2;
mem[16'hAB3D] = 8'hD6;
mem[16'hAB3E] = 8'hBF;
mem[16'hAB3F] = 8'hCC;
mem[16'hAB40] = 8'hD3;
mem[16'hAB41] = 8'hCD;
mem[16'hAB42] = 8'hC9;
mem[16'hAB43] = 8'hBC;
mem[16'hAB44] = 8'hD4;
mem[16'hAB45] = 8'hCE;
mem[16'hAB46] = 8'hCA;
mem[16'hAB47] = 8'hBD;
mem[16'hAB48] = 8'hD5;
mem[16'hAB49] = 8'hCF;
mem[16'hAB4A] = 8'hCB;
mem[16'hAB4B] = 8'hBE;
mem[16'hAB4C] = 8'hD6;
mem[16'hAB4D] = 8'hD2;
mem[16'hAB4E] = 8'hCC;
mem[16'hAB4F] = 8'hBF;
mem[16'hAB50] = 8'hD7;
mem[16'hAB51] = 8'hDC;
mem[16'hAB52] = 8'hE4;
mem[16'hAB53] = 8'hE9;
mem[16'hAB54] = 8'hD9;
mem[16'hAB55] = 8'hDD;
mem[16'hAB56] = 8'hE5;
mem[16'hAB57] = 8'hEA;
mem[16'hAB58] = 8'hDA;
mem[16'hAB59] = 8'hDE;
mem[16'hAB5A] = 8'hE6;
mem[16'hAB5B] = 8'hEB;
mem[16'hAB5C] = 8'hDB;
mem[16'hAB5D] = 8'hDF;
mem[16'hAB5E] = 8'hE7;
mem[16'hAB5F] = 8'hEC;
mem[16'hAB60] = 8'hFF;
mem[16'hAB61] = 8'h4C;
mem[16'hAB62] = 8'h73;
mem[16'hAB63] = 8'hB3;
mem[16'hAB64] = 8'hA9;
mem[16'hAB65] = 8'h00;
mem[16'hAB66] = 8'h9D;
mem[16'hAB67] = 8'hE8;
mem[16'hAB68] = 8'hB4;
mem[16'hAB69] = 8'hA9;
mem[16'hAB6A] = 8'h01;
mem[16'hAB6B] = 8'h9D;
mem[16'hAB6C] = 8'hE7;
mem[16'hAB6D] = 8'hB4;
mem[16'hAB6E] = 8'h8E;
mem[16'hAB6F] = 8'h9C;
mem[16'hAB70] = 8'hB3;
mem[16'hAB71] = 8'h20;
mem[16'hAB72] = 8'h44;
mem[16'hAB73] = 8'hB2;
mem[16'hAB74] = 8'hAE;
mem[16'hAB75] = 8'h9C;
mem[16'hAB76] = 8'hB3;
mem[16'hAB77] = 8'h9D;
mem[16'hAB78] = 8'hC7;
mem[16'hAB79] = 8'hB4;
mem[16'hAB7A] = 8'h8D;
mem[16'hAB7B] = 8'hD2;
mem[16'hAB7C] = 8'hB5;
mem[16'hAB7D] = 8'h8D;
mem[16'hAB7E] = 8'hD4;
mem[16'hAB7F] = 8'hB5;
mem[16'hAB80] = 8'hAD;
mem[16'hAB81] = 8'hF1;
mem[16'hAB82] = 8'hB5;
mem[16'hAB83] = 8'h9D;
mem[16'hAB84] = 8'hC6;
mem[16'hAB85] = 8'hB4;
mem[16'hAB86] = 8'h8D;
mem[16'hAB87] = 8'hD1;
mem[16'hAB88] = 8'hB5;
mem[16'hAB89] = 8'h8D;
mem[16'hAB8A] = 8'hD3;
mem[16'hAB8B] = 8'hB5;
mem[16'hAB8C] = 8'hAD;
mem[16'hAB8D] = 8'hC2;
mem[16'hAB8E] = 8'hB5;
mem[16'hAB8F] = 8'h9D;
mem[16'hAB90] = 8'hC8;
mem[16'hAB91] = 8'hB4;
mem[16'hAB92] = 8'h20;
mem[16'hAB93] = 8'h37;
mem[16'hAB94] = 8'hB0;
mem[16'hAB95] = 8'h20;
mem[16'hAB96] = 8'h0C;
mem[16'hAB97] = 8'hAF;
mem[16'hAB98] = 8'h20;
mem[16'hAB99] = 8'hD6;
mem[16'hAB9A] = 8'hB7;
mem[16'hAB9B] = 8'h20;
mem[16'hAB9C] = 8'h3A;
mem[16'hAB9D] = 8'hAF;
mem[16'hAB9E] = 8'hAE;
mem[16'hAB9F] = 8'h9C;
mem[16'hABA0] = 8'hB3;
mem[16'hABA1] = 8'hA9;
mem[16'hABA2] = 8'h06;
mem[16'hABA3] = 8'h8D;
mem[16'hABA4] = 8'hC5;
mem[16'hABA5] = 8'hB5;
mem[16'hABA6] = 8'hBD;
mem[16'hABA7] = 8'hC6;
mem[16'hABA8] = 8'hB4;
mem[16'hABA9] = 8'h8D;
mem[16'hABAA] = 8'hD1;
mem[16'hABAB] = 8'hB5;
mem[16'hABAC] = 8'hBD;
mem[16'hABAD] = 8'hC7;
mem[16'hABAE] = 8'hB4;
mem[16'hABAF] = 8'h8D;
mem[16'hABB0] = 8'hD2;
mem[16'hABB1] = 8'hB5;
mem[16'hABB2] = 8'hBD;
mem[16'hABB3] = 8'hC8;
mem[16'hABB4] = 8'hB4;
mem[16'hABB5] = 8'h8D;
mem[16'hABB6] = 8'hC2;
mem[16'hABB7] = 8'hB5;
mem[16'hABB8] = 8'h8D;
mem[16'hABB9] = 8'hF6;
mem[16'hABBA] = 8'hB5;
mem[16'hABBB] = 8'hBD;
mem[16'hABBC] = 8'hE7;
mem[16'hABBD] = 8'hB4;
mem[16'hABBE] = 8'h8D;
mem[16'hABBF] = 8'hEE;
mem[16'hABC0] = 8'hB5;
mem[16'hABC1] = 8'hBD;
mem[16'hABC2] = 8'hE8;
mem[16'hABC3] = 8'hB4;
mem[16'hABC4] = 8'h8D;
mem[16'hABC5] = 8'hEF;
mem[16'hABC6] = 8'hB5;
mem[16'hABC7] = 8'h8E;
mem[16'hABC8] = 8'hD9;
mem[16'hABC9] = 8'hB5;
mem[16'hABCA] = 8'hA9;
mem[16'hABCB] = 8'hFF;
mem[16'hABCC] = 8'h8D;
mem[16'hABCD] = 8'hE0;
mem[16'hABCE] = 8'hB5;
mem[16'hABCF] = 8'h8D;
mem[16'hABD0] = 8'hE1;
mem[16'hABD1] = 8'hB5;
mem[16'hABD2] = 8'hAD;
mem[16'hABD3] = 8'hE2;
mem[16'hABD4] = 8'hB3;
mem[16'hABD5] = 8'h8D;
mem[16'hABD6] = 8'hDA;
mem[16'hABD7] = 8'hB5;
mem[16'hABD8] = 8'h18;
mem[16'hABD9] = 8'h4C;
mem[16'hABDA] = 8'h5E;
mem[16'hABDB] = 8'hAF;
mem[16'hABDC] = 8'hA9;
mem[16'hABDD] = 8'h00;
mem[16'hABDE] = 8'hAA;
mem[16'hABDF] = 8'h9D;
mem[16'hABE0] = 8'hD1;
mem[16'hABE1] = 8'hB5;
mem[16'hABE2] = 8'hE8;
mem[16'hABE3] = 8'hE0;
mem[16'hABE4] = 8'h2D;
mem[16'hABE5] = 8'hD0;
mem[16'hABE6] = 8'hF8;
mem[16'hABE7] = 8'hAD;
mem[16'hABE8] = 8'hBF;
mem[16'hABE9] = 8'hB5;
mem[16'hABEA] = 8'h49;
mem[16'hABEB] = 8'hFF;
mem[16'hABEC] = 8'h8D;
mem[16'hABED] = 8'hF9;
mem[16'hABEE] = 8'hB5;
mem[16'hABEF] = 8'hAD;
mem[16'hABF0] = 8'hC0;
mem[16'hABF1] = 8'hB5;
mem[16'hABF2] = 8'h8D;
mem[16'hABF3] = 8'hF8;
mem[16'hABF4] = 8'hB5;
mem[16'hABF5] = 8'hAD;
mem[16'hABF6] = 8'hC1;
mem[16'hABF7] = 8'hB5;
mem[16'hABF8] = 8'h0A;
mem[16'hABF9] = 8'h0A;
mem[16'hABFA] = 8'h0A;
mem[16'hABFB] = 8'h0A;
mem[16'hABFC] = 8'hAA;
mem[16'hABFD] = 8'h8E;
mem[16'hABFE] = 8'hF7;
mem[16'hABFF] = 8'hB5;
mem[16'hAC00] = 8'h05;
mem[16'hAC01] = 8'h07;
mem[16'hAC02] = 8'h05;
mem[16'hAC03] = 8'h03;
mem[16'hAC04] = 8'h05;
mem[16'hAC05] = 8'h07;
mem[16'hAC06] = 8'h05;
mem[16'hAC07] = 8'h19;
mem[16'hAC08] = 8'h17;
mem[16'hAC09] = 8'h11;
mem[16'hAC0A] = 8'h13;
mem[16'hAC0B] = 8'h11;
mem[16'hAC0C] = 8'h17;
mem[16'hAC0D] = 8'h18;
mem[16'hAC0E] = 8'h18;
mem[16'hAC0F] = 8'h18;
mem[16'hAC10] = 8'h00;
mem[16'hAC11] = 8'h00;
mem[16'hAC12] = 8'h00;
mem[16'hAC13] = 8'h00;
mem[16'hAC14] = 8'h71;
mem[16'hAC15] = 8'h73;
mem[16'hAC16] = 8'h71;
mem[16'hAC17] = 8'h77;
mem[16'hAC18] = 8'h79;
mem[16'hAC19] = 8'h7B;
mem[16'hAC1A] = 8'h79;
mem[16'hAC1B] = 8'h65;
mem[16'hAC1C] = 8'h63;
mem[16'hAC1D] = 8'h65;
mem[16'hAC1E] = 8'h67;
mem[16'hAC1F] = 8'h65;
mem[16'hAC20] = 8'h5B;
mem[16'hAC21] = 8'h54;
mem[16'hAC22] = 8'h54;
mem[16'hAC23] = 8'h54;
mem[16'hAC24] = 8'h54;
mem[16'hAC25] = 8'h54;
mem[16'hAC26] = 8'h54;
mem[16'hAC27] = 8'h54;
mem[16'hAC28] = 8'h60;
mem[16'hAC29] = 8'h60;
mem[16'hAC2A] = 8'h60;
mem[16'hAC2B] = 8'h60;
mem[16'hAC2C] = 8'h69;
mem[16'hAC2D] = 8'h6B;
mem[16'hAC2E] = 8'h69;
mem[16'hAC2F] = 8'h6F;
mem[16'hAC30] = 8'h71;
mem[16'hAC31] = 8'h73;
mem[16'hAC32] = 8'h71;
mem[16'hAC33] = 8'h6D;
mem[16'hAC34] = 8'h6B;
mem[16'hAC35] = 8'h6D;
mem[16'hAC36] = 8'h6F;
mem[16'hAC37] = 8'h6D;
mem[16'hAC38] = 8'h63;
mem[16'hAC39] = 8'h6C;
mem[16'hAC3A] = 8'h6C;
mem[16'hAC3B] = 8'h6C;
mem[16'hAC3C] = 8'h6C;
mem[16'hAC3D] = 8'h6C;
mem[16'hAC3E] = 8'h6C;
mem[16'hAC3F] = 8'h6C;
mem[16'hAC40] = 8'hDC;
mem[16'hAC41] = 8'hC6;
mem[16'hAC42] = 8'h43;
mem[16'hAC43] = 8'h52;
mem[16'hAC44] = 8'h5D;
mem[16'hAC45] = 8'h6C;
mem[16'hAC46] = 8'hA8;
mem[16'hAC47] = 8'h46;
mem[16'hAC48] = 8'h5A;
mem[16'hAC49] = 8'h50;
mem[16'hAC4A] = 8'h63;
mem[16'hAC4B] = 8'hA4;
mem[16'hAC4C] = 8'h4E;
mem[16'hAC4D] = 8'h7D;
mem[16'hAC4E] = 8'h51;
mem[16'hAC4F] = 8'hC3;
mem[16'hAC50] = 8'hE0;
mem[16'hAC51] = 8'h4F;
mem[16'hAC52] = 8'hDE;
mem[16'hAC53] = 8'hC8;
mem[16'hAC54] = 8'h48;
mem[16'hAC55] = 8'hB5;
mem[16'hAC56] = 8'h85;
mem[16'hAC57] = 8'h48;
mem[16'hAC58] = 8'h59;
mem[16'hAC59] = 8'h49;
mem[16'hAC5A] = 8'h43;
mem[16'hAC5B] = 8'h3E;
mem[16'hAC5C] = 8'hF5;
mem[16'hAC5D] = 8'h41;
mem[16'hAC5E] = 8'hF9;
mem[16'hAC5F] = 8'hF9;
mem[16'hAC60] = 8'h66;
mem[16'hAC61] = 8'h70;
mem[16'hAC62] = 8'h28;
mem[16'hAC63] = 8'h65;
mem[16'hAC64] = 8'h80;
mem[16'hAC65] = 8'h74;
mem[16'hAC66] = 8'h2F;
mem[16'hAC67] = 8'h61;
mem[16'hAC68] = 8'h8C;
mem[16'hAC69] = 8'hA5;
mem[16'hAC6A] = 8'h8A;
mem[16'hAC6B] = 8'hA0;
mem[16'hAC6C] = 8'h73;
mem[16'hAC6D] = 8'h8D;
mem[16'hAC6E] = 8'hB9;
mem[16'hAC6F] = 8'h70;
mem[16'hAC70] = 8'h71;
mem[16'hAC71] = 8'h2B;
mem[16'hAC72] = 8'h6B;
mem[16'hAC73] = 8'hEF;
mem[16'hAC74] = 8'h20;
mem[16'hAC75] = 8'h74;
mem[16'hAC76] = 8'h66;
mem[16'hAC77] = 8'h6E;
mem[16'hAC78] = 8'h1D;
mem[16'hAC79] = 8'hD0;
mem[16'hAC7A] = 8'h66;
mem[16'hAC7B] = 8'h39;
mem[16'hAC7C] = 8'hDA;
mem[16'hAC7D] = 8'h7B;
mem[16'hAC7E] = 8'h6F;
mem[16'hAC7F] = 8'h21;
mem[16'hAC80] = 8'h86;
mem[16'hAC81] = 8'h65;
mem[16'hAC82] = 8'h93;
mem[16'hAC83] = 8'hDE;
mem[16'hAC84] = 8'h82;
mem[16'hAC85] = 8'h61;
mem[16'hAC86] = 8'h4A;
mem[16'hAC87] = 8'h0B;
mem[16'hAC88] = 8'h24;
mem[16'hAC89] = 8'h96;
mem[16'hAC8A] = 8'h06;
mem[16'hAC8B] = 8'h8F;
mem[16'hAC8C] = 8'h8C;
mem[16'hAC8D] = 8'hAC;
mem[16'hAC8E] = 8'hE1;
mem[16'hAC8F] = 8'h96;
mem[16'hAC90] = 8'h70;
mem[16'hAC91] = 8'h42;
mem[16'hAC92] = 8'h8D;
mem[16'hAC93] = 8'h1F;
mem[16'hAC94] = 8'h38;
mem[16'hAC95] = 8'h8A;
mem[16'hAC96] = 8'h1A;
mem[16'hAC97] = 8'h8E;
mem[16'hAC98] = 8'h85;
mem[16'hAC99] = 8'h15;
mem[16'hAC9A] = 8'h9E;
mem[16'hAC9B] = 8'h9B;
mem[16'hAC9C] = 8'h78;
mem[16'hAC9D] = 8'h11;
mem[16'hAC9E] = 8'h90;
mem[16'hAC9F] = 8'h82;
mem[16'hACA0] = 8'hAC;
mem[16'hACA1] = 8'h0D;
mem[16'hACA2] = 8'h66;
mem[16'hACA3] = 8'h9E;
mem[16'hACA4] = 8'h4A;
mem[16'hACA5] = 8'h45;
mem[16'hACA6] = 8'h9C;
mem[16'hACA7] = 8'hA7;
mem[16'hACA8] = 8'h24;
mem[16'hACA9] = 8'h05;
mem[16'hACAA] = 8'h07;
mem[16'hACAB] = 8'h05;
mem[16'hACAC] = 8'h03;
mem[16'hACAD] = 8'h05;
mem[16'hACAE] = 8'h07;
mem[16'hACAF] = 8'h05;
mem[16'hACB0] = 8'h3C;
mem[16'hACB1] = 8'h46;
mem[16'hACB2] = 8'h19;
mem[16'hACB3] = 8'h17;
mem[16'hACB4] = 8'h11;
mem[16'hACB5] = 8'h13;
mem[16'hACB6] = 8'h11;
mem[16'hACB7] = 8'h17;
mem[16'hACB8] = 8'h58;
mem[16'hACB9] = 8'h18;
mem[16'hACBA] = 8'h18;
mem[16'hACBB] = 8'h18;
mem[16'hACBC] = 8'h00;
mem[16'hACBD] = 8'h00;
mem[16'hACBE] = 8'h00;
mem[16'hACBF] = 8'h00;
mem[16'hACC0] = 8'hD9;
mem[16'hACC1] = 8'h4D;
mem[16'hACC2] = 8'hB4;
mem[16'hACC3] = 8'hC3;
mem[16'hACC4] = 8'h24;
mem[16'hACC5] = 8'h16;
mem[16'hACC6] = 8'hD9;
mem[16'hACC7] = 8'h4B;
mem[16'hACC8] = 8'h64;
mem[16'hACC9] = 8'h71;
mem[16'hACCA] = 8'h73;
mem[16'hACCB] = 8'h71;
mem[16'hACCC] = 8'h77;
mem[16'hACCD] = 8'h79;
mem[16'hACCE] = 8'h7B;
mem[16'hACCF] = 8'h79;
mem[16'hACD0] = 8'h3E;
mem[16'hACD1] = 8'h5D;
mem[16'hACD2] = 8'h65;
mem[16'hACD3] = 8'h63;
mem[16'hACD4] = 8'h65;
mem[16'hACD5] = 8'h67;
mem[16'hACD6] = 8'h65;
mem[16'hACD7] = 8'h5B;
mem[16'hACD8] = 8'hBE;
mem[16'hACD9] = 8'h54;
mem[16'hACDA] = 8'h54;
mem[16'hACDB] = 8'h54;
mem[16'hACDC] = 8'h54;
mem[16'hACDD] = 8'h54;
mem[16'hACDE] = 8'h54;
mem[16'hACDF] = 8'h54;
mem[16'hACE0] = 8'h0E;
mem[16'hACE1] = 8'hE4;
mem[16'hACE2] = 8'h0E;
mem[16'hACE3] = 8'h42;
mem[16'hACE4] = 8'h60;
mem[16'hACE5] = 8'h60;
mem[16'hACE6] = 8'h60;
mem[16'hACE7] = 8'h60;
mem[16'hACE8] = 8'hF1;
mem[16'hACE9] = 8'h69;
mem[16'hACEA] = 8'h6B;
mem[16'hACEB] = 8'h69;
mem[16'hACEC] = 8'h6F;
mem[16'hACED] = 8'h71;
mem[16'hACEE] = 8'h73;
mem[16'hACEF] = 8'h71;
mem[16'hACF0] = 8'hDC;
mem[16'hACF1] = 8'hD0;
mem[16'hACF2] = 8'h6D;
mem[16'hACF3] = 8'h6B;
mem[16'hACF4] = 8'h6D;
mem[16'hACF5] = 8'h6F;
mem[16'hACF6] = 8'h6D;
mem[16'hACF7] = 8'h63;
mem[16'hACF8] = 8'hD9;
mem[16'hACF9] = 8'h6C;
mem[16'hACFA] = 8'h6C;
mem[16'hACFB] = 8'h6C;
mem[16'hACFC] = 8'h6C;
mem[16'hACFD] = 8'h6C;
mem[16'hACFE] = 8'h6C;
mem[16'hACFF] = 8'h6C;
mem[16'hAD00] = 8'hB3;
mem[16'hAD01] = 8'hBD;
mem[16'hAD02] = 8'hC8;
mem[16'hAD03] = 8'hB4;
mem[16'hAD04] = 8'h29;
mem[16'hAD05] = 8'h7F;
mem[16'hAD06] = 8'h0D;
mem[16'hAD07] = 8'h9E;
mem[16'hAD08] = 8'hB3;
mem[16'hAD09] = 8'h9D;
mem[16'hAD0A] = 8'hC8;
mem[16'hAD0B] = 8'hB4;
mem[16'hAD0C] = 8'h20;
mem[16'hAD0D] = 8'h37;
mem[16'hAD0E] = 8'hB0;
mem[16'hAD0F] = 8'h4C;
mem[16'hAD10] = 8'h7F;
mem[16'hAD11] = 8'hB3;
mem[16'hAD12] = 8'h20;
mem[16'hAD13] = 8'h00;
mem[16'hAD14] = 8'hB3;
mem[16'hAD15] = 8'h4C;
mem[16'hAD16] = 8'h7F;
mem[16'hAD17] = 8'hB3;
mem[16'hAD18] = 8'h20;
mem[16'hAD19] = 8'h28;
mem[16'hAD1A] = 8'hAB;
mem[16'hAD1B] = 8'h20;
mem[16'hAD1C] = 8'hB6;
mem[16'hAD1D] = 8'hB0;
mem[16'hAD1E] = 8'hB0;
mem[16'hAD1F] = 8'hEF;
mem[16'hAD20] = 8'hEE;
mem[16'hAD21] = 8'hE4;
mem[16'hAD22] = 8'hB5;
mem[16'hAD23] = 8'hD0;
mem[16'hAD24] = 8'hF6;
mem[16'hAD25] = 8'hEE;
mem[16'hAD26] = 8'hE5;
mem[16'hAD27] = 8'hB5;
mem[16'hAD28] = 8'h4C;
mem[16'hAD29] = 8'h1B;
mem[16'hAD2A] = 8'hAD;
mem[16'hAD2B] = 8'h20;
mem[16'hAD2C] = 8'h28;
mem[16'hAD2D] = 8'hAB;
mem[16'hAD2E] = 8'hAE;
mem[16'hAD2F] = 8'h9C;
mem[16'hAD30] = 8'hB3;
mem[16'hAD31] = 8'hBD;
mem[16'hAD32] = 8'hC8;
mem[16'hAD33] = 8'hB4;
mem[16'hAD34] = 8'h10;
mem[16'hAD35] = 8'h03;
mem[16'hAD36] = 8'h4C;
mem[16'hAD37] = 8'h7B;
mem[16'hAD38] = 8'hB3;
mem[16'hAD39] = 8'hAE;
mem[16'hAD3A] = 8'h9C;
mem[16'hAD3B] = 8'hB3;
mem[16'hAD3C] = 8'hBD;
mem[16'hAD3D] = 8'hC6;
mem[16'hAD3E] = 8'hB4;
mem[16'hAD3F] = 8'h8D;
mem[16'hAD40] = 8'hD1;
mem[16'hAD41] = 8'hB5;
mem[16'hAD42] = 8'h9D;
mem[16'hAD43] = 8'hE6;
mem[16'hAD44] = 8'hB4;
mem[16'hAD45] = 8'hA9;
mem[16'hAD46] = 8'hFF;
mem[16'hAD47] = 8'h9D;
mem[16'hAD48] = 8'hC6;
mem[16'hAD49] = 8'hB4;
mem[16'hAD4A] = 8'hBC;
mem[16'hAD4B] = 8'hC7;
mem[16'hAD4C] = 8'hB4;
mem[16'hAD4D] = 8'h8C;
mem[16'hAD4E] = 8'hD2;
mem[16'hAD4F] = 8'hB5;
mem[16'hAD50] = 8'h20;
mem[16'hAD51] = 8'h37;
mem[16'hAD52] = 8'hB0;
mem[16'hAD53] = 8'h18;
mem[16'hAD54] = 8'h20;
mem[16'hAD55] = 8'h5E;
mem[16'hAD56] = 8'hAF;
mem[16'hAD57] = 8'hB0;
mem[16'hAD58] = 8'h2A;
mem[16'hAD59] = 8'h20;
mem[16'hAD5A] = 8'h0C;
mem[16'hAD5B] = 8'hAF;
mem[16'hAD5C] = 8'hA0;
mem[16'hAD5D] = 8'h0C;
mem[16'hAD5E] = 8'h8C;
mem[16'hAD5F] = 8'h9C;
mem[16'hAD60] = 8'hB3;
mem[16'hAD61] = 8'hB1;
mem[16'hAD62] = 8'h42;
mem[16'hAD63] = 8'h30;
mem[16'hAD64] = 8'h0B;
mem[16'hAD65] = 8'hF0;
mem[16'hAD66] = 8'h09;
mem[16'hAD67] = 8'h48;
mem[16'hAD68] = 8'hC8;
mem[16'hAD69] = 8'hB1;
mem[16'hAD6A] = 8'h42;
mem[16'hAD6B] = 8'hA8;
mem[16'hAD6C] = 8'h68;
mem[16'hAD6D] = 8'h20;
mem[16'hAD6E] = 8'h89;
mem[16'hAD6F] = 8'hAD;
mem[16'hAD70] = 8'hAC;
mem[16'hAD71] = 8'h9C;
mem[16'hAD72] = 8'hB3;
mem[16'hAD73] = 8'hC8;
mem[16'hAD74] = 8'hC8;
mem[16'hAD75] = 8'hD0;
mem[16'hAD76] = 8'hE7;
mem[16'hAD77] = 8'hAD;
mem[16'hAD78] = 8'hD3;
mem[16'hAD79] = 8'hB5;
mem[16'hAD7A] = 8'hAC;
mem[16'hAD7B] = 8'hD4;
mem[16'hAD7C] = 8'hB5;
mem[16'hAD7D] = 8'h20;
mem[16'hAD7E] = 8'h89;
mem[16'hAD7F] = 8'hAD;
mem[16'hAD80] = 8'h38;
mem[16'hAD81] = 8'hB0;
mem[16'hAD82] = 8'hD1;
mem[16'hAD83] = 8'h20;
mem[16'hAD84] = 8'hFB;
mem[16'hAD85] = 8'hAF;
mem[16'hAD86] = 8'h4C;
mem[16'hAD87] = 8'h7F;
mem[16'hAD88] = 8'hB3;
mem[16'hAD89] = 8'h38;
mem[16'hAD8A] = 8'h20;
mem[16'hAD8B] = 8'hDD;
mem[16'hAD8C] = 8'hB2;
mem[16'hAD8D] = 8'hA9;
mem[16'hAD8E] = 8'h00;
mem[16'hAD8F] = 8'hA2;
mem[16'hAD90] = 8'h05;
mem[16'hAD91] = 8'h9D;
mem[16'hAD92] = 8'hF0;
mem[16'hAD93] = 8'hB5;
mem[16'hAD94] = 8'hCA;
mem[16'hAD95] = 8'h10;
mem[16'hAD96] = 8'hFA;
mem[16'hAD97] = 8'h60;
mem[16'hAD98] = 8'h20;
mem[16'hAD99] = 8'hDC;
mem[16'hAD9A] = 8'hAB;
mem[16'hAD9B] = 8'hA9;
mem[16'hAD9C] = 8'hFF;
mem[16'hAD9D] = 8'h8D;
mem[16'hAD9E] = 8'hF9;
mem[16'hAD9F] = 8'hB5;
mem[16'hADA0] = 8'h20;
mem[16'hADA1] = 8'hF7;
mem[16'hADA2] = 8'hAF;
mem[16'hADA3] = 8'hA9;
mem[16'hADA4] = 8'h16;
mem[16'hADA5] = 8'h8D;
mem[16'hADA6] = 8'h9D;
mem[16'hADA7] = 8'hB3;
mem[16'hADA8] = 8'h20;
mem[16'hADA9] = 8'h00;
mem[16'hADAA] = 8'h00;
mem[16'hADAB] = 8'h00;
mem[16'hADAC] = 8'h00;
mem[16'hADAD] = 8'h00;
mem[16'hADAE] = 8'h00;
mem[16'hADAF] = 8'h00;
mem[16'hADB0] = 8'hBD;
mem[16'hADB1] = 8'hAF;
mem[16'hADB2] = 8'h00;
mem[16'hADB3] = 8'h00;
mem[16'hADB4] = 8'h00;
mem[16'hADB5] = 8'h00;
mem[16'hADB6] = 8'h00;
mem[16'hADB7] = 8'h00;
mem[16'hADB8] = 8'hF7;
mem[16'hADB9] = 8'h00;
mem[16'hADBA] = 8'h00;
mem[16'hADBB] = 8'h00;
mem[16'hADBC] = 8'h40;
mem[16'hADBD] = 8'h40;
mem[16'hADBE] = 8'h40;
mem[16'hADBF] = 8'h40;
mem[16'hADC0] = 8'h20;
mem[16'hADC1] = 8'h42;
mem[16'hADC2] = 8'hAE;
mem[16'hADC3] = 8'h20;
mem[16'hADC4] = 8'h2F;
mem[16'hADC5] = 8'hAE;
mem[16'hADC6] = 8'h20;
mem[16'hADC7] = 8'h2F;
mem[16'hADC8] = 8'hAE;
mem[16'hADC9] = 8'h40;
mem[16'hADCA] = 8'h40;
mem[16'hADCB] = 8'h40;
mem[16'hADCC] = 8'h40;
mem[16'hADCD] = 8'h40;
mem[16'hADCE] = 8'h40;
mem[16'hADCF] = 8'h40;
mem[16'hADD0] = 8'h00;
mem[16'hADD1] = 8'h8E;
mem[16'hADD2] = 8'h40;
mem[16'hADD3] = 8'h40;
mem[16'hADD4] = 8'h40;
mem[16'hADD5] = 8'h40;
mem[16'hADD6] = 8'h40;
mem[16'hADD7] = 8'h80;
mem[16'hADD8] = 8'h53;
mem[16'hADD9] = 8'h80;
mem[16'hADDA] = 8'h80;
mem[16'hADDB] = 8'h80;
mem[16'hADDC] = 8'h80;
mem[16'hADDD] = 8'h80;
mem[16'hADDE] = 8'h80;
mem[16'hADDF] = 8'h80;
mem[16'hADE0] = 8'h10;
mem[16'hADE1] = 8'h02;
mem[16'hADE2] = 8'hA0;
mem[16'hADE3] = 8'hAA;
mem[16'hADE4] = 8'h80;
mem[16'hADE5] = 8'h80;
mem[16'hADE6] = 8'h80;
mem[16'hADE7] = 8'h80;
mem[16'hADE8] = 8'hBD;
mem[16'hADE9] = 8'h80;
mem[16'hADEA] = 8'h80;
mem[16'hADEB] = 8'h80;
mem[16'hADEC] = 8'h80;
mem[16'hADED] = 8'hC0;
mem[16'hADEE] = 8'hC0;
mem[16'hADEF] = 8'hC0;
mem[16'hADF0] = 8'h0A;
mem[16'hADF1] = 8'hB0;
mem[16'hADF2] = 8'hC0;
mem[16'hADF3] = 8'hC0;
mem[16'hADF4] = 8'hC0;
mem[16'hADF5] = 8'hC0;
mem[16'hADF6] = 8'hC0;
mem[16'hADF7] = 8'hC0;
mem[16'hADF8] = 8'hB3;
mem[16'hADF9] = 8'hC0;
mem[16'hADFA] = 8'hC0;
mem[16'hADFB] = 8'hC0;
mem[16'hADFC] = 8'hC0;
mem[16'hADFD] = 8'hC0;
mem[16'hADFE] = 8'hC0;
mem[16'hADFF] = 8'hC0;
mem[16'hAE00] = 8'hFD;
mem[16'hAE01] = 8'hBD;
mem[16'hAE02] = 8'hE7;
mem[16'hAE03] = 8'hB4;
mem[16'hAE04] = 8'h85;
mem[16'hAE05] = 8'h44;
mem[16'hAE06] = 8'hBD;
mem[16'hAE07] = 8'hE8;
mem[16'hAE08] = 8'hB4;
mem[16'hAE09] = 8'h85;
mem[16'hAE0A] = 8'h45;
mem[16'hAE0B] = 8'h20;
mem[16'hAE0C] = 8'h42;
mem[16'hAE0D] = 8'hAE;
mem[16'hAE0E] = 8'hA9;
mem[16'hAE0F] = 8'hA0;
mem[16'hAE10] = 8'h20;
mem[16'hAE11] = 8'hED;
mem[16'hAE12] = 8'hFD;
mem[16'hAE13] = 8'hE8;
mem[16'hAE14] = 8'hE8;
mem[16'hAE15] = 8'hE8;
mem[16'hAE16] = 8'hA0;
mem[16'hAE17] = 8'h1D;
mem[16'hAE18] = 8'hBD;
mem[16'hAE19] = 8'hC6;
mem[16'hAE1A] = 8'hB4;
mem[16'hAE1B] = 8'h20;
mem[16'hAE1C] = 8'hED;
mem[16'hAE1D] = 8'hFD;
mem[16'hAE1E] = 8'hE8;
mem[16'hAE1F] = 8'h88;
mem[16'hAE20] = 8'h10;
mem[16'hAE21] = 8'hF6;
mem[16'hAE22] = 8'h20;
mem[16'hAE23] = 8'h2F;
mem[16'hAE24] = 8'hAE;
mem[16'hAE25] = 8'h20;
mem[16'hAE26] = 8'h30;
mem[16'hAE27] = 8'hB2;
mem[16'hAE28] = 8'h90;
mem[16'hAE29] = 8'hA7;
mem[16'hAE2A] = 8'hB0;
mem[16'hAE2B] = 8'h9E;
mem[16'hAE2C] = 8'h4C;
mem[16'hAE2D] = 8'h7F;
mem[16'hAE2E] = 8'hB3;
mem[16'hAE2F] = 8'hA9;
mem[16'hAE30] = 8'h8D;
mem[16'hAE31] = 8'h20;
mem[16'hAE32] = 8'hED;
mem[16'hAE33] = 8'hFD;
mem[16'hAE34] = 8'hCE;
mem[16'hAE35] = 8'h9D;
mem[16'hAE36] = 8'hB3;
mem[16'hAE37] = 8'hD0;
mem[16'hAE38] = 8'h08;
mem[16'hAE39] = 8'h20;
mem[16'hAE3A] = 8'h0C;
mem[16'hAE3B] = 8'hFD;
mem[16'hAE3C] = 8'hA9;
mem[16'hAE3D] = 8'h15;
mem[16'hAE3E] = 8'h8D;
mem[16'hAE3F] = 8'h9D;
mem[16'hAE40] = 8'hB3;
mem[16'hAE41] = 8'h60;
mem[16'hAE42] = 8'hA0;
mem[16'hAE43] = 8'h02;
mem[16'hAE44] = 8'hA9;
mem[16'hAE45] = 8'h00;
mem[16'hAE46] = 8'h48;
mem[16'hAE47] = 8'hA5;
mem[16'hAE48] = 8'h44;
mem[16'hAE49] = 8'hD9;
mem[16'hAE4A] = 8'hA4;
mem[16'hAE4B] = 8'hB3;
mem[16'hAE4C] = 8'h90;
mem[16'hAE4D] = 8'h12;
mem[16'hAE4E] = 8'hF9;
mem[16'hAE4F] = 8'hA4;
mem[16'hAE50] = 8'hB3;
mem[16'hAE51] = 8'h85;
mem[16'hAE52] = 8'h44;
mem[16'hAE53] = 8'hA5;
mem[16'hAE54] = 8'h45;
mem[16'hAE55] = 8'hE9;
mem[16'hAE56] = 8'h00;
mem[16'hAE57] = 8'h85;
mem[16'hAE58] = 8'h45;
mem[16'hAE59] = 8'h68;
mem[16'hAE5A] = 8'h69;
mem[16'hAE5B] = 8'h00;
mem[16'hAE5C] = 8'h48;
mem[16'hAE5D] = 8'h4C;
mem[16'hAE5E] = 8'h47;
mem[16'hAE5F] = 8'hAE;
mem[16'hAE60] = 8'h68;
mem[16'hAE61] = 8'h09;
mem[16'hAE62] = 8'hB0;
mem[16'hAE63] = 8'h20;
mem[16'hAE64] = 8'hED;
mem[16'hAE65] = 8'hFD;
mem[16'hAE66] = 8'h88;
mem[16'hAE67] = 8'h10;
mem[16'hAE68] = 8'hDB;
mem[16'hAE69] = 8'h60;
mem[16'hAE6A] = 8'h20;
mem[16'hAE6B] = 8'h08;
mem[16'hAE6C] = 8'hAF;
mem[16'hAE6D] = 8'hA0;
mem[16'hAE6E] = 8'h00;
mem[16'hAE6F] = 8'h8C;
mem[16'hAE70] = 8'hC5;
mem[16'hAE71] = 8'hB5;
mem[16'hAE72] = 8'hB1;
mem[16'hAE73] = 8'h42;
mem[16'hAE74] = 8'h99;
mem[16'hAE75] = 8'hD1;
mem[16'hAE76] = 8'hB5;
mem[16'hAE77] = 8'hC8;
mem[16'hAE78] = 8'hC0;
mem[16'hAE79] = 8'h2D;
mem[16'hAE7A] = 8'hD0;
mem[16'hAE7B] = 8'hF6;
mem[16'hAE7C] = 8'h18;
mem[16'hAE7D] = 8'h60;
mem[16'hAE7E] = 8'h20;
mem[16'hAE7F] = 8'h08;
mem[16'hAE80] = 8'hAF;
mem[16'hAE81] = 8'hA0;
mem[16'hAE82] = 8'h00;
mem[16'hAE83] = 8'hB9;
mem[16'hAE84] = 8'hD1;
mem[16'hAE85] = 8'hB5;
mem[16'hAE86] = 8'h91;
mem[16'hAE87] = 8'h42;
mem[16'hAE88] = 8'hC8;
mem[16'hAE89] = 8'hC0;
mem[16'hAE8A] = 8'h2D;
mem[16'hAE8B] = 8'hD0;
mem[16'hAE8C] = 8'hF6;
mem[16'hAE8D] = 8'h60;
mem[16'hAE8E] = 8'h20;
mem[16'hAE8F] = 8'hDC;
mem[16'hAE90] = 8'hAB;
mem[16'hAE91] = 8'hA9;
mem[16'hAE92] = 8'h04;
mem[16'hAE93] = 8'h20;
mem[16'hAE94] = 8'h58;
mem[16'hAE95] = 8'hB0;
mem[16'hAE96] = 8'hAD;
mem[16'hAE97] = 8'hF9;
mem[16'hAE98] = 8'hB5;
mem[16'hAE99] = 8'h49;
mem[16'hAE9A] = 8'hFF;
mem[16'hAE9B] = 8'h8D;
mem[16'hAE9C] = 8'hC1;
mem[16'hAE9D] = 8'hB3;
mem[16'hAE9E] = 8'hA9;
mem[16'hAE9F] = 8'h11;
mem[16'hAEA0] = 8'h8D;
mem[16'hAEA1] = 8'hEB;
mem[16'hAEA2] = 8'hB3;
mem[16'hAEA3] = 8'hA9;
mem[16'hAEA4] = 8'h01;
mem[16'hAEA5] = 8'h8D;
mem[16'hAEA6] = 8'hEC;
mem[16'hAEA7] = 8'hB3;
mem[16'hAEA8] = 8'hA2;
mem[16'hAEA9] = 8'h00;
mem[16'hAEAA] = 8'h01;
mem[16'hAEAB] = 8'h02;
mem[16'hAEAC] = 8'h03;
mem[16'hAEAD] = 8'h04;
mem[16'hAEAE] = 8'h05;
mem[16'hAEAF] = 8'h06;
mem[16'hAEB0] = 8'hD0;
mem[16'hAEB1] = 8'hFA;
mem[16'hAEB2] = 8'h07;
mem[16'hAEB3] = 8'h08;
mem[16'hAEB4] = 8'h09;
mem[16'hAEB5] = 8'h0A;
mem[16'hAEB6] = 8'h0B;
mem[16'hAEB7] = 8'h0C;
mem[16'hAEB8] = 8'hA0;
mem[16'hAEB9] = 8'h0D;
mem[16'hAEBA] = 8'h0E;
mem[16'hAEBB] = 8'h0F;
mem[16'hAEBC] = 8'h00;
mem[16'hAEBD] = 8'h01;
mem[16'hAEBE] = 8'h02;
mem[16'hAEBF] = 8'h03;
mem[16'hAEC0] = 8'hE8;
mem[16'hAEC1] = 8'h88;
mem[16'hAEC2] = 8'h10;
mem[16'hAEC3] = 8'hF6;
mem[16'hAEC4] = 8'hE0;
mem[16'hAEC5] = 8'h44;
mem[16'hAEC6] = 8'hD0;
mem[16'hAEC7] = 8'hEC;
mem[16'hAEC8] = 8'hA2;
mem[16'hAEC9] = 8'h04;
mem[16'hAECA] = 8'h05;
mem[16'hAECB] = 8'h06;
mem[16'hAECC] = 8'h07;
mem[16'hAECD] = 8'h08;
mem[16'hAECE] = 8'h09;
mem[16'hAECF] = 8'h0A;
mem[16'hAED0] = 8'h00;
mem[16'hAED1] = 8'h8A;
mem[16'hAED2] = 8'h0B;
mem[16'hAED3] = 8'h0C;
mem[16'hAED4] = 8'h0D;
mem[16'hAED5] = 8'h0E;
mem[16'hAED6] = 8'h0F;
mem[16'hAED7] = 8'h00;
mem[16'hAED8] = 8'h20;
mem[16'hAED9] = 8'h01;
mem[16'hAEDA] = 8'h02;
mem[16'hAEDB] = 8'h03;
mem[16'hAEDC] = 8'h04;
mem[16'hAEDD] = 8'h05;
mem[16'hAEDE] = 8'h06;
mem[16'hAEDF] = 8'h07;
mem[16'hAEE0] = 8'h88;
mem[16'hAEE1] = 8'h88;
mem[16'hAEE2] = 8'h8D;
mem[16'hAEE3] = 8'hEC;
mem[16'hAEE4] = 8'h08;
mem[16'hAEE5] = 8'h09;
mem[16'hAEE6] = 8'h0A;
mem[16'hAEE7] = 8'h0B;
mem[16'hAEE8] = 8'h8C;
mem[16'hAEE9] = 8'h0C;
mem[16'hAEEA] = 8'h0D;
mem[16'hAEEB] = 8'h0E;
mem[16'hAEEC] = 8'h0F;
mem[16'hAEED] = 8'h00;
mem[16'hAEEE] = 8'h01;
mem[16'hAEEF] = 8'h02;
mem[16'hAEF0] = 8'h02;
mem[16'hAEF1] = 8'h20;
mem[16'hAEF2] = 8'h03;
mem[16'hAEF3] = 8'h04;
mem[16'hAEF4] = 8'h05;
mem[16'hAEF5] = 8'h06;
mem[16'hAEF6] = 8'h07;
mem[16'hAEF7] = 8'h08;
mem[16'hAEF8] = 8'h30;
mem[16'hAEF9] = 8'h09;
mem[16'hAEFA] = 8'h0A;
mem[16'hAEFB] = 8'h0B;
mem[16'hAEFC] = 8'h0C;
mem[16'hAEFD] = 8'h0D;
mem[16'hAEFE] = 8'h0E;
mem[16'hAEFF] = 8'h0F;
mem[16'hAF00] = 8'hC2;
mem[16'hAF01] = 8'hB7;
mem[16'hAF02] = 8'h20;
mem[16'hAF03] = 8'h4A;
mem[16'hAF04] = 8'hB7;
mem[16'hAF05] = 8'h4C;
mem[16'hAF06] = 8'h7F;
mem[16'hAF07] = 8'hB3;
mem[16'hAF08] = 8'hA2;
mem[16'hAF09] = 8'h00;
mem[16'hAF0A] = 8'hF0;
mem[16'hAF0B] = 8'h06;
mem[16'hAF0C] = 8'hA2;
mem[16'hAF0D] = 8'h02;
mem[16'hAF0E] = 8'hD0;
mem[16'hAF0F] = 8'h02;
mem[16'hAF10] = 8'hA2;
mem[16'hAF11] = 8'h04;
mem[16'hAF12] = 8'hBD;
mem[16'hAF13] = 8'hC7;
mem[16'hAF14] = 8'hB5;
mem[16'hAF15] = 8'h85;
mem[16'hAF16] = 8'h42;
mem[16'hAF17] = 8'hBD;
mem[16'hAF18] = 8'hC8;
mem[16'hAF19] = 8'hB5;
mem[16'hAF1A] = 8'h85;
mem[16'hAF1B] = 8'h43;
mem[16'hAF1C] = 8'h60;
mem[16'hAF1D] = 8'h2C;
mem[16'hAF1E] = 8'hD5;
mem[16'hAF1F] = 8'hB5;
mem[16'hAF20] = 8'h70;
mem[16'hAF21] = 8'h01;
mem[16'hAF22] = 8'h60;
mem[16'hAF23] = 8'h20;
mem[16'hAF24] = 8'hE4;
mem[16'hAF25] = 8'hAF;
mem[16'hAF26] = 8'hA9;
mem[16'hAF27] = 8'h02;
mem[16'hAF28] = 8'h20;
mem[16'hAF29] = 8'h52;
mem[16'hAF2A] = 8'hB0;
mem[16'hAF2B] = 8'hA9;
mem[16'hAF2C] = 8'hBF;
mem[16'hAF2D] = 8'h2D;
mem[16'hAF2E] = 8'hD5;
mem[16'hAF2F] = 8'hB5;
mem[16'hAF30] = 8'h8D;
mem[16'hAF31] = 8'hD5;
mem[16'hAF32] = 8'hB5;
mem[16'hAF33] = 8'h60;
mem[16'hAF34] = 8'hAD;
mem[16'hAF35] = 8'hD5;
mem[16'hAF36] = 8'hB5;
mem[16'hAF37] = 8'h30;
mem[16'hAF38] = 8'h01;
mem[16'hAF39] = 8'h60;
mem[16'hAF3A] = 8'h20;
mem[16'hAF3B] = 8'h4B;
mem[16'hAF3C] = 8'hAF;
mem[16'hAF3D] = 8'hA9;
mem[16'hAF3E] = 8'h02;
mem[16'hAF3F] = 8'h20;
mem[16'hAF40] = 8'h52;
mem[16'hAF41] = 8'hB0;
mem[16'hAF42] = 8'hA9;
mem[16'hAF43] = 8'h7F;
mem[16'hAF44] = 8'h2D;
mem[16'hAF45] = 8'hD5;
mem[16'hAF46] = 8'hB5;
mem[16'hAF47] = 8'h8D;
mem[16'hAF48] = 8'hD5;
mem[16'hAF49] = 8'hB5;
mem[16'hAF4A] = 8'h60;
mem[16'hAF4B] = 8'hAD;
mem[16'hAF4C] = 8'hC9;
mem[16'hAF4D] = 8'hB5;
mem[16'hAF4E] = 8'h8D;
mem[16'hAF4F] = 8'hF0;
mem[16'hAF50] = 8'hB7;
mem[16'hAF51] = 8'hAD;
mem[16'hAF52] = 8'hCA;
mem[16'hAF53] = 8'hB5;
mem[16'hAF54] = 8'h8D;
mem[16'hAF55] = 8'hF1;
mem[16'hAF56] = 8'hB7;
mem[16'hAF57] = 8'hAE;
mem[16'hAF58] = 8'hD3;
mem[16'hAF59] = 8'hB5;
mem[16'hAF5A] = 8'hAC;
mem[16'hAF5B] = 8'hD4;
mem[16'hAF5C] = 8'hB5;
mem[16'hAF5D] = 8'h60;
mem[16'hAF5E] = 8'h08;
mem[16'hAF5F] = 8'h20;
mem[16'hAF60] = 8'h34;
mem[16'hAF61] = 8'hAF;
mem[16'hAF62] = 8'h20;
mem[16'hAF63] = 8'h4B;
mem[16'hAF64] = 8'hAF;
mem[16'hAF65] = 8'h20;
mem[16'hAF66] = 8'h0C;
mem[16'hAF67] = 8'hAF;
mem[16'hAF68] = 8'h28;
mem[16'hAF69] = 8'hB0;
mem[16'hAF6A] = 8'h09;
mem[16'hAF6B] = 8'hAE;
mem[16'hAF6C] = 8'hD1;
mem[16'hAF6D] = 8'hB5;
mem[16'hAF6E] = 8'hAC;
mem[16'hAF6F] = 8'hD2;
mem[16'hAF70] = 8'hB5;
mem[16'hAF71] = 8'h4C;
mem[16'hAF72] = 8'hB5;
mem[16'hAF73] = 8'hAF;
mem[16'hAF74] = 8'hA0;
mem[16'hAF75] = 8'h01;
mem[16'hAF76] = 8'hB1;
mem[16'hAF77] = 8'h42;
mem[16'hAF78] = 8'hF0;
mem[16'hAF79] = 8'h08;
mem[16'hAF7A] = 8'hAA;
mem[16'hAF7B] = 8'hC8;
mem[16'hAF7C] = 8'hB1;
mem[16'hAF7D] = 8'h42;
mem[16'hAF7E] = 8'hA8;
mem[16'hAF7F] = 8'h4C;
mem[16'hAF80] = 8'hB5;
mem[16'hAF81] = 8'hAF;
mem[16'hAF82] = 8'hAD;
mem[16'hAF83] = 8'hBB;
mem[16'hAF84] = 8'hB5;
mem[16'hAF85] = 8'hC9;
mem[16'hAF86] = 8'h04;
mem[16'hAF87] = 8'hF0;
mem[16'hAF88] = 8'h02;
mem[16'hAF89] = 8'h38;
mem[16'hAF8A] = 8'h60;
mem[16'hAF8B] = 8'h20;
mem[16'hAF8C] = 8'h44;
mem[16'hAF8D] = 8'hB2;
mem[16'hAF8E] = 8'hA0;
mem[16'hAF8F] = 8'h02;
mem[16'hAF90] = 8'h91;
mem[16'hAF91] = 8'h42;
mem[16'hAF92] = 8'h48;
mem[16'hAF93] = 8'h88;
mem[16'hAF94] = 8'hAD;
mem[16'hAF95] = 8'hF1;
mem[16'hAF96] = 8'hB5;
mem[16'hAF97] = 8'h91;
mem[16'hAF98] = 8'h42;
mem[16'hAF99] = 8'h48;
mem[16'hAF9A] = 8'h20;
mem[16'hAF9B] = 8'h3A;
mem[16'hAF9C] = 8'hAF;
mem[16'hAF9D] = 8'h20;
mem[16'hAF9E] = 8'hD6;
mem[16'hAF9F] = 8'hB7;
mem[16'hAFA0] = 8'hA0;
mem[16'hAFA1] = 8'h05;
mem[16'hAFA2] = 8'hAD;
mem[16'hAFA3] = 8'hDE;
mem[16'hAFA4] = 8'hB5;
mem[16'hAFA5] = 8'h91;
mem[16'hAFA6] = 8'h42;
mem[16'hAFA7] = 8'hC8;
mem[16'hAFA8] = 8'hAD;
mem[16'hAFA9] = 8'h00;
mem[16'hAFAA] = 8'h00;
mem[16'hAFAB] = 8'h00;
mem[16'hAFAC] = 8'h00;
mem[16'hAFAD] = 8'h10;
mem[16'hAFAE] = 8'h10;
mem[16'hAFAF] = 8'h10;
mem[16'hAFB0] = 8'hA8;
mem[16'hAFB1] = 8'hA9;
mem[16'hAFB2] = 8'h10;
mem[16'hAFB3] = 8'h20;
mem[16'hAFB4] = 8'h20;
mem[16'hAFB5] = 8'h20;
mem[16'hAFB6] = 8'h20;
mem[16'hAFB7] = 8'h30;
mem[16'hAFB8] = 8'hD3;
mem[16'hAFB9] = 8'h30;
mem[16'hAFBA] = 8'h30;
mem[16'hAFBB] = 8'h30;
mem[16'hAFBC] = 8'h40;
mem[16'hAFBD] = 8'h40;
mem[16'hAFBE] = 8'h40;
mem[16'hAFBF] = 8'h40;
mem[16'hAFC0] = 8'hA0;
mem[16'hAFC1] = 8'h05;
mem[16'hAFC2] = 8'hB1;
mem[16'hAFC3] = 8'h42;
mem[16'hAFC4] = 8'h8D;
mem[16'hAFC5] = 8'hDC;
mem[16'hAFC6] = 8'hB5;
mem[16'hAFC7] = 8'h18;
mem[16'hAFC8] = 8'h6D;
mem[16'hAFC9] = 8'h50;
mem[16'hAFCA] = 8'h50;
mem[16'hAFCB] = 8'h50;
mem[16'hAFCC] = 8'h50;
mem[16'hAFCD] = 8'h60;
mem[16'hAFCE] = 8'h60;
mem[16'hAFCF] = 8'h60;
mem[16'hAFD0] = 8'h42;
mem[16'hAFD1] = 8'h8D;
mem[16'hAFD2] = 8'h60;
mem[16'hAFD3] = 8'h70;
mem[16'hAFD4] = 8'h70;
mem[16'hAFD5] = 8'h70;
mem[16'hAFD6] = 8'h70;
mem[16'hAFD7] = 8'h80;
mem[16'hAFD8] = 8'hDF;
mem[16'hAFD9] = 8'h80;
mem[16'hAFDA] = 8'h80;
mem[16'hAFDB] = 8'h80;
mem[16'hAFDC] = 8'h90;
mem[16'hAFDD] = 8'h90;
mem[16'hAFDE] = 8'h90;
mem[16'hAFDF] = 8'h90;
mem[16'hAFE0] = 8'h01;
mem[16'hAFE1] = 8'h4C;
mem[16'hAFE2] = 8'h52;
mem[16'hAFE3] = 8'hB0;
mem[16'hAFE4] = 8'hA0;
mem[16'hAFE5] = 8'hA0;
mem[16'hAFE6] = 8'hA0;
mem[16'hAFE7] = 8'hA0;
mem[16'hAFE8] = 8'hCC;
mem[16'hAFE9] = 8'hB0;
mem[16'hAFEA] = 8'hB0;
mem[16'hAFEB] = 8'hB0;
mem[16'hAFEC] = 8'hB0;
mem[16'hAFED] = 8'hC0;
mem[16'hAFEE] = 8'hC0;
mem[16'hAFEF] = 8'hC0;
mem[16'hAFF0] = 8'hAE;
mem[16'hAFF1] = 8'hD6;
mem[16'hAFF2] = 8'hC0;
mem[16'hAFF3] = 8'hD0;
mem[16'hAFF4] = 8'hD0;
mem[16'hAFF5] = 8'hD0;
mem[16'hAFF6] = 8'hD0;
mem[16'hAFF7] = 8'hE0;
mem[16'hAFF8] = 8'h01;
mem[16'hAFF9] = 8'hE0;
mem[16'hAFFA] = 8'hE0;
mem[16'hAFFB] = 8'hE0;
mem[16'hAFFC] = 8'hF0;
mem[16'hAFFD] = 8'hF0;
mem[16'hAFFE] = 8'hF0;
mem[16'hAFFF] = 8'hF0;
mem[16'hB000] = 8'h8C;
mem[16'hB001] = 8'hF0;
mem[16'hB002] = 8'hB7;
mem[16'hB003] = 8'hAC;
mem[16'hB004] = 8'hC4;
mem[16'hB005] = 8'hAA;
mem[16'hB006] = 8'h8C;
mem[16'hB007] = 8'hF1;
mem[16'hB008] = 8'hB7;
mem[16'hB009] = 8'hAE;
mem[16'hB00A] = 8'hFA;
mem[16'hB00B] = 8'hB5;
mem[16'hB00C] = 8'hA0;
mem[16'hB00D] = 8'h00;
mem[16'hB00E] = 8'h4C;
mem[16'hB00F] = 8'h52;
mem[16'hB010] = 8'hB0;
mem[16'hB011] = 8'h08;
mem[16'hB012] = 8'h20;
mem[16'hB013] = 8'h45;
mem[16'hB014] = 8'hB0;
mem[16'hB015] = 8'h28;
mem[16'hB016] = 8'hB0;
mem[16'hB017] = 8'h08;
mem[16'hB018] = 8'hAC;
mem[16'hB019] = 8'hBD;
mem[16'hB01A] = 8'hB3;
mem[16'hB01B] = 8'hAE;
mem[16'hB01C] = 8'hBC;
mem[16'hB01D] = 8'hB3;
mem[16'hB01E] = 8'hD0;
mem[16'hB01F] = 8'h0A;
mem[16'hB020] = 8'hAE;
mem[16'hB021] = 8'hBC;
mem[16'hB022] = 8'hB4;
mem[16'hB023] = 8'hD0;
mem[16'hB024] = 8'h02;
mem[16'hB025] = 8'h38;
mem[16'hB026] = 8'h60;
mem[16'hB027] = 8'hAC;
mem[16'hB028] = 8'hBD;
mem[16'hB029] = 8'hB4;
mem[16'hB02A] = 8'h8E;
mem[16'hB02B] = 8'h97;
mem[16'hB02C] = 8'hB3;
mem[16'hB02D] = 8'h8C;
mem[16'hB02E] = 8'h98;
mem[16'hB02F] = 8'hB3;
mem[16'hB030] = 8'hA9;
mem[16'hB031] = 8'h01;
mem[16'hB032] = 8'h20;
mem[16'hB033] = 8'h52;
mem[16'hB034] = 8'hB0;
mem[16'hB035] = 8'h18;
mem[16'hB036] = 8'h60;
mem[16'hB037] = 8'h20;
mem[16'hB038] = 8'h45;
mem[16'hB039] = 8'hB0;
mem[16'hB03A] = 8'hAE;
mem[16'hB03B] = 8'h97;
mem[16'hB03C] = 8'hB3;
mem[16'hB03D] = 8'hAC;
mem[16'hB03E] = 8'h98;
mem[16'hB03F] = 8'hB3;
mem[16'hB040] = 8'hA9;
mem[16'hB041] = 8'h02;
mem[16'hB042] = 8'h4C;
mem[16'hB043] = 8'h52;
mem[16'hB044] = 8'hB0;
mem[16'hB045] = 8'hAD;
mem[16'hB046] = 8'hC5;
mem[16'hB047] = 8'hAA;
mem[16'hB048] = 8'h8D;
mem[16'hB049] = 8'hF0;
mem[16'hB04A] = 8'hB7;
mem[16'hB04B] = 8'hAD;
mem[16'hB04C] = 8'hC6;
mem[16'hB04D] = 8'hAA;
mem[16'hB04E] = 8'h8D;
mem[16'hB04F] = 8'hF1;
mem[16'hB050] = 8'hB7;
mem[16'hB051] = 8'h60;
mem[16'hB052] = 8'h8E;
mem[16'hB053] = 8'hEC;
mem[16'hB054] = 8'hB7;
mem[16'hB055] = 8'h8C;
mem[16'hB056] = 8'hED;
mem[16'hB057] = 8'hB7;
mem[16'hB058] = 8'h8D;
mem[16'hB059] = 8'hF4;
mem[16'hB05A] = 8'hB7;
mem[16'hB05B] = 8'hC9;
mem[16'hB05C] = 8'h02;
mem[16'hB05D] = 8'hD0;
mem[16'hB05E] = 8'h06;
mem[16'hB05F] = 8'h0D;
mem[16'hB060] = 8'hD5;
mem[16'hB061] = 8'hB5;
mem[16'hB062] = 8'h8D;
mem[16'hB063] = 8'hD5;
mem[16'hB064] = 8'hB5;
mem[16'hB065] = 8'hAD;
mem[16'hB066] = 8'hF9;
mem[16'hB067] = 8'hB5;
mem[16'hB068] = 8'h49;
mem[16'hB069] = 8'hFF;
mem[16'hB06A] = 8'h8D;
mem[16'hB06B] = 8'hEB;
mem[16'hB06C] = 8'hB7;
mem[16'hB06D] = 8'hAD;
mem[16'hB06E] = 8'hF7;
mem[16'hB06F] = 8'hB5;
mem[16'hB070] = 8'h8D;
mem[16'hB071] = 8'hE9;
mem[16'hB072] = 8'hB7;
mem[16'hB073] = 8'hAD;
mem[16'hB074] = 8'hF8;
mem[16'hB075] = 8'hB5;
mem[16'hB076] = 8'h8D;
mem[16'hB077] = 8'hEA;
mem[16'hB078] = 8'hB7;
mem[16'hB079] = 8'hAD;
mem[16'hB07A] = 8'hE2;
mem[16'hB07B] = 8'hB5;
mem[16'hB07C] = 8'h8D;
mem[16'hB07D] = 8'hF2;
mem[16'hB07E] = 8'hB7;
mem[16'hB07F] = 8'hAD;
mem[16'hB080] = 8'hE3;
mem[16'hB081] = 8'hB5;
mem[16'hB082] = 8'h8D;
mem[16'hB083] = 8'hF3;
mem[16'hB084] = 8'hB7;
mem[16'hB085] = 8'hA9;
mem[16'hB086] = 8'h01;
mem[16'hB087] = 8'h8D;
mem[16'hB088] = 8'hE8;
mem[16'hB089] = 8'hB7;
mem[16'hB08A] = 8'hAC;
mem[16'hB08B] = 8'hC1;
mem[16'hB08C] = 8'hAA;
mem[16'hB08D] = 8'hAD;
mem[16'hB08E] = 8'hC2;
mem[16'hB08F] = 8'hAA;
mem[16'hB090] = 8'h20;
mem[16'hB091] = 8'hB5;
mem[16'hB092] = 8'hB7;
mem[16'hB093] = 8'hAD;
mem[16'hB094] = 8'hF6;
mem[16'hB095] = 8'hB7;
mem[16'hB096] = 8'h8D;
mem[16'hB097] = 8'hBF;
mem[16'hB098] = 8'hB5;
mem[16'hB099] = 8'hA9;
mem[16'hB09A] = 8'hFF;
mem[16'hB09B] = 8'h8D;
mem[16'hB09C] = 8'hEB;
mem[16'hB09D] = 8'hB7;
mem[16'hB09E] = 8'hB0;
mem[16'hB09F] = 8'h01;
mem[16'hB0A0] = 8'h60;
mem[16'hB0A1] = 8'hAD;
mem[16'hB0A2] = 8'hF5;
mem[16'hB0A3] = 8'hB7;
mem[16'hB0A4] = 8'hA0;
mem[16'hB0A5] = 8'h07;
mem[16'hB0A6] = 8'hC9;
mem[16'hB0A7] = 8'h20;
mem[16'hB0A8] = 8'hF0;
mem[16'hB0A9] = 8'h00;
mem[16'hB0AA] = 8'h01;
mem[16'hB0AB] = 8'h02;
mem[16'hB0AC] = 8'h03;
mem[16'hB0AD] = 8'h00;
mem[16'hB0AE] = 8'h01;
mem[16'hB0AF] = 8'h02;
mem[16'hB0B0] = 8'hA0;
mem[16'hB0B1] = 8'h08;
mem[16'hB0B2] = 8'h03;
mem[16'hB0B3] = 8'h00;
mem[16'hB0B4] = 8'h01;
mem[16'hB0B5] = 8'h02;
mem[16'hB0B6] = 8'h03;
mem[16'hB0B7] = 8'h00;
mem[16'hB0B8] = 8'hB5;
mem[16'hB0B9] = 8'h01;
mem[16'hB0BA] = 8'h02;
mem[16'hB0BB] = 8'h03;
mem[16'hB0BC] = 8'h00;
mem[16'hB0BD] = 8'h01;
mem[16'hB0BE] = 8'h02;
mem[16'hB0BF] = 8'h03;
mem[16'hB0C0] = 8'hB5;
mem[16'hB0C1] = 8'hCD;
mem[16'hB0C2] = 8'hE1;
mem[16'hB0C3] = 8'hB5;
mem[16'hB0C4] = 8'hF0;
mem[16'hB0C5] = 8'h66;
mem[16'hB0C6] = 8'h20;
mem[16'hB0C7] = 8'h1D;
mem[16'hB0C8] = 8'hAF;
mem[16'hB0C9] = 8'h00;
mem[16'hB0CA] = 8'h01;
mem[16'hB0CB] = 8'h02;
mem[16'hB0CC] = 8'h03;
mem[16'hB0CD] = 8'h00;
mem[16'hB0CE] = 8'h01;
mem[16'hB0CF] = 8'h02;
mem[16'hB0D0] = 8'h1C;
mem[16'hB0D1] = 8'hD0;
mem[16'hB0D2] = 8'h03;
mem[16'hB0D3] = 8'h00;
mem[16'hB0D4] = 8'h01;
mem[16'hB0D5] = 8'h02;
mem[16'hB0D6] = 8'h03;
mem[16'hB0D7] = 8'h00;
mem[16'hB0D8] = 8'hB5;
mem[16'hB0D9] = 8'h01;
mem[16'hB0DA] = 8'h02;
mem[16'hB0DB] = 8'h03;
mem[16'hB0DC] = 8'h00;
mem[16'hB0DD] = 8'h01;
mem[16'hB0DE] = 8'h02;
mem[16'hB0DF] = 8'h03;
mem[16'hB0E0] = 8'hB5;
mem[16'hB0E1] = 8'h90;
mem[16'hB0E2] = 8'h10;
mem[16'hB0E3] = 8'hD0;
mem[16'hB0E4] = 8'h00;
mem[16'hB0E5] = 8'h01;
mem[16'hB0E6] = 8'h02;
mem[16'hB0E7] = 8'h03;
mem[16'hB0E8] = 8'hCD;
mem[16'hB0E9] = 8'h00;
mem[16'hB0EA] = 8'h01;
mem[16'hB0EB] = 8'h02;
mem[16'hB0EC] = 8'h03;
mem[16'hB0ED] = 8'h00;
mem[16'hB0EE] = 8'h01;
mem[16'hB0EF] = 8'h02;
mem[16'hB0F0] = 8'h90;
mem[16'hB0F1] = 8'hD7;
mem[16'hB0F2] = 8'h03;
mem[16'hB0F3] = 8'h00;
mem[16'hB0F4] = 8'h01;
mem[16'hB0F5] = 8'h02;
mem[16'hB0F6] = 8'h03;
mem[16'hB0F7] = 8'h00;
mem[16'hB0F8] = 8'hDC;
mem[16'hB0F9] = 8'h01;
mem[16'hB0FA] = 8'h02;
mem[16'hB0FB] = 8'h03;
mem[16'hB0FC] = 8'h00;
mem[16'hB0FD] = 8'h01;
mem[16'hB0FE] = 8'h02;
mem[16'hB0FF] = 8'h03;
mem[16'hB100] = 8'hAF;
mem[16'hB101] = 8'hB1;
mem[16'hB102] = 8'h42;
mem[16'hB103] = 8'hD0;
mem[16'hB104] = 8'h0F;
mem[16'hB105] = 8'hAD;
mem[16'hB106] = 8'hBB;
mem[16'hB107] = 8'hB5;
mem[16'hB108] = 8'hC9;
mem[16'hB109] = 8'h04;
mem[16'hB10A] = 8'hF0;
mem[16'hB10B] = 8'h02;
mem[16'hB10C] = 8'h38;
mem[16'hB10D] = 8'h60;
mem[16'hB10E] = 8'h20;
mem[16'hB10F] = 8'h34;
mem[16'hB110] = 8'hB1;
mem[16'hB111] = 8'h4C;
mem[16'hB112] = 8'h20;
mem[16'hB113] = 8'hB1;
mem[16'hB114] = 8'h8D;
mem[16'hB115] = 8'hD6;
mem[16'hB116] = 8'hB5;
mem[16'hB117] = 8'hC8;
mem[16'hB118] = 8'hB1;
mem[16'hB119] = 8'h42;
mem[16'hB11A] = 8'h8D;
mem[16'hB11B] = 8'hD7;
mem[16'hB11C] = 8'hB5;
mem[16'hB11D] = 8'h20;
mem[16'hB11E] = 8'hDC;
mem[16'hB11F] = 8'hAF;
mem[16'hB120] = 8'hAD;
mem[16'hB121] = 8'hE4;
mem[16'hB122] = 8'hB5;
mem[16'hB123] = 8'h8D;
mem[16'hB124] = 8'hE0;
mem[16'hB125] = 8'hB5;
mem[16'hB126] = 8'hAD;
mem[16'hB127] = 8'hE5;
mem[16'hB128] = 8'hB5;
mem[16'hB129] = 8'h8D;
mem[16'hB12A] = 8'hE1;
mem[16'hB12B] = 8'hB5;
mem[16'hB12C] = 8'h20;
mem[16'hB12D] = 8'h10;
mem[16'hB12E] = 8'hAF;
mem[16'hB12F] = 8'hAC;
mem[16'hB130] = 8'hE6;
mem[16'hB131] = 8'hB5;
mem[16'hB132] = 8'h18;
mem[16'hB133] = 8'h60;
mem[16'hB134] = 8'h8C;
mem[16'hB135] = 8'h9D;
mem[16'hB136] = 8'hB3;
mem[16'hB137] = 8'h20;
mem[16'hB138] = 8'h44;
mem[16'hB139] = 8'hB2;
mem[16'hB13A] = 8'hAC;
mem[16'hB13B] = 8'h9D;
mem[16'hB13C] = 8'hB3;
mem[16'hB13D] = 8'hC8;
mem[16'hB13E] = 8'h91;
mem[16'hB13F] = 8'h42;
mem[16'hB140] = 8'h8D;
mem[16'hB141] = 8'hD7;
mem[16'hB142] = 8'hB5;
mem[16'hB143] = 8'h88;
mem[16'hB144] = 8'hAD;
mem[16'hB145] = 8'hF1;
mem[16'hB146] = 8'hB5;
mem[16'hB147] = 8'h91;
mem[16'hB148] = 8'h42;
mem[16'hB149] = 8'h8D;
mem[16'hB14A] = 8'hD6;
mem[16'hB14B] = 8'hB5;
mem[16'hB14C] = 8'h20;
mem[16'hB14D] = 8'h10;
mem[16'hB14E] = 8'hAF;
mem[16'hB14F] = 8'h20;
mem[16'hB150] = 8'hD6;
mem[16'hB151] = 8'hB7;
mem[16'hB152] = 8'hA9;
mem[16'hB153] = 8'hC0;
mem[16'hB154] = 8'h0D;
mem[16'hB155] = 8'hD5;
mem[16'hB156] = 8'hB5;
mem[16'hB157] = 8'h8D;
mem[16'hB158] = 8'hD5;
mem[16'hB159] = 8'hB5;
mem[16'hB15A] = 8'h60;
mem[16'hB15B] = 8'hAE;
mem[16'hB15C] = 8'hEA;
mem[16'hB15D] = 8'hB5;
mem[16'hB15E] = 8'h8E;
mem[16'hB15F] = 8'hBD;
mem[16'hB160] = 8'hB5;
mem[16'hB161] = 8'hAE;
mem[16'hB162] = 8'hEB;
mem[16'hB163] = 8'hB5;
mem[16'hB164] = 8'h8E;
mem[16'hB165] = 8'hBE;
mem[16'hB166] = 8'hB5;
mem[16'hB167] = 8'hAE;
mem[16'hB168] = 8'hEC;
mem[16'hB169] = 8'hB5;
mem[16'hB16A] = 8'hAC;
mem[16'hB16B] = 8'hED;
mem[16'hB16C] = 8'hB5;
mem[16'hB16D] = 8'h8E;
mem[16'hB16E] = 8'hBF;
mem[16'hB16F] = 8'hB5;
mem[16'hB170] = 8'h8C;
mem[16'hB171] = 8'hC0;
mem[16'hB172] = 8'hB5;
mem[16'hB173] = 8'hE8;
mem[16'hB174] = 8'hD0;
mem[16'hB175] = 8'h01;
mem[16'hB176] = 8'hC8;
mem[16'hB177] = 8'hCC;
mem[16'hB178] = 8'hE9;
mem[16'hB179] = 8'hB5;
mem[16'hB17A] = 8'hD0;
mem[16'hB17B] = 8'h11;
mem[16'hB17C] = 8'hEC;
mem[16'hB17D] = 8'hE8;
mem[16'hB17E] = 8'hB5;
mem[16'hB17F] = 8'hD0;
mem[16'hB180] = 8'h0C;
mem[16'hB181] = 8'hA2;
mem[16'hB182] = 8'h00;
mem[16'hB183] = 8'hA0;
mem[16'hB184] = 8'h00;
mem[16'hB185] = 8'hEE;
mem[16'hB186] = 8'hEA;
mem[16'hB187] = 8'hB5;
mem[16'hB188] = 8'hD0;
mem[16'hB189] = 8'h03;
mem[16'hB18A] = 8'hEE;
mem[16'hB18B] = 8'hEB;
mem[16'hB18C] = 8'hB5;
mem[16'hB18D] = 8'h8E;
mem[16'hB18E] = 8'hEC;
mem[16'hB18F] = 8'hB5;
mem[16'hB190] = 8'h8C;
mem[16'hB191] = 8'hED;
mem[16'hB192] = 8'hB5;
mem[16'hB193] = 8'h60;
mem[16'hB194] = 8'hEE;
mem[16'hB195] = 8'hE6;
mem[16'hB196] = 8'hB5;
mem[16'hB197] = 8'hD0;
mem[16'hB198] = 8'h08;
mem[16'hB199] = 8'hEE;
mem[16'hB19A] = 8'hE4;
mem[16'hB19B] = 8'hB5;
mem[16'hB19C] = 8'hD0;
mem[16'hB19D] = 8'h03;
mem[16'hB19E] = 8'hEE;
mem[16'hB19F] = 8'hE5;
mem[16'hB1A0] = 8'hB5;
mem[16'hB1A1] = 8'h60;
mem[16'hB1A2] = 8'hAC;
mem[16'hB1A3] = 8'hC3;
mem[16'hB1A4] = 8'hB5;
mem[16'hB1A5] = 8'hAE;
mem[16'hB1A6] = 8'hC4;
mem[16'hB1A7] = 8'hB5;
mem[16'hB1A8] = 8'h84;
mem[16'hB1A9] = 8'h00;
mem[16'hB1AA] = 8'h04;
mem[16'hB1AB] = 8'h08;
mem[16'hB1AC] = 8'h0C;
mem[16'hB1AD] = 8'h10;
mem[16'hB1AE] = 8'h14;
mem[16'hB1AF] = 8'h18;
mem[16'hB1B0] = 8'h03;
mem[16'hB1B1] = 8'hEE;
mem[16'hB1B2] = 8'h1C;
mem[16'hB1B3] = 8'h20;
mem[16'hB1B4] = 8'h24;
mem[16'hB1B5] = 8'h28;
mem[16'hB1B6] = 8'h2C;
mem[16'hB1B7] = 8'h30;
mem[16'hB1B8] = 8'hD0;
mem[16'hB1B9] = 8'h34;
mem[16'hB1BA] = 8'h38;
mem[16'hB1BB] = 8'h3C;
mem[16'hB1BC] = 8'h40;
mem[16'hB1BD] = 8'h44;
mem[16'hB1BE] = 8'h48;
mem[16'hB1BF] = 8'h4C;
mem[16'hB1C0] = 8'hC2;
mem[16'hB1C1] = 8'hB5;
mem[16'hB1C2] = 8'hCE;
mem[16'hB1C3] = 8'hC1;
mem[16'hB1C4] = 8'hB5;
mem[16'hB1C5] = 8'h60;
mem[16'hB1C6] = 8'h4C;
mem[16'hB1C7] = 8'h7F;
mem[16'hB1C8] = 8'hB3;
mem[16'hB1C9] = 8'h50;
mem[16'hB1CA] = 8'h54;
mem[16'hB1CB] = 8'h58;
mem[16'hB1CC] = 8'h5C;
mem[16'hB1CD] = 8'h60;
mem[16'hB1CE] = 8'h64;
mem[16'hB1CF] = 8'h68;
mem[16'hB1D0] = 8'h42;
mem[16'hB1D1] = 8'hAD;
mem[16'hB1D2] = 8'h6C;
mem[16'hB1D3] = 8'h70;
mem[16'hB1D4] = 8'h74;
mem[16'hB1D5] = 8'h78;
mem[16'hB1D6] = 8'h7C;
mem[16'hB1D7] = 8'h80;
mem[16'hB1D8] = 8'h8D;
mem[16'hB1D9] = 8'h84;
mem[16'hB1DA] = 8'h88;
mem[16'hB1DB] = 8'h8C;
mem[16'hB1DC] = 8'h90;
mem[16'hB1DD] = 8'h94;
mem[16'hB1DE] = 8'h98;
mem[16'hB1DF] = 8'h9C;
mem[16'hB1E0] = 8'h18;
mem[16'hB1E1] = 8'hEE;
mem[16'hB1E2] = 8'hD8;
mem[16'hB1E3] = 8'hB5;
mem[16'hB1E4] = 8'hA0;
mem[16'hB1E5] = 8'hA4;
mem[16'hB1E6] = 8'hA8;
mem[16'hB1E7] = 8'hAC;
mem[16'hB1E8] = 8'h51;
mem[16'hB1E9] = 8'hB0;
mem[16'hB1EA] = 8'hB4;
mem[16'hB1EB] = 8'hB8;
mem[16'hB1EC] = 8'hBC;
mem[16'hB1ED] = 8'hC0;
mem[16'hB1EE] = 8'hC4;
mem[16'hB1EF] = 8'hC8;
mem[16'hB1F0] = 8'hB4;
mem[16'hB1F1] = 8'hF0;
mem[16'hB1F2] = 8'hCC;
mem[16'hB1F3] = 8'hD0;
mem[16'hB1F4] = 8'hD4;
mem[16'hB1F5] = 8'hD8;
mem[16'hB1F6] = 8'hDC;
mem[16'hB1F7] = 8'hE0;
mem[16'hB1F8] = 8'hE8;
mem[16'hB1F9] = 8'hE4;
mem[16'hB1FA] = 8'hE8;
mem[16'hB1FB] = 8'hEC;
mem[16'hB1FC] = 8'hF0;
mem[16'hB1FD] = 8'hF4;
mem[16'hB1FE] = 8'hF8;
mem[16'hB1FF] = 8'hFC;
mem[16'hB200] = 8'h8C;
mem[16'hB201] = 8'hED;
mem[16'hB202] = 8'hAE;
mem[16'hB203] = 8'hAF;
mem[16'hB204] = 8'hA8;
mem[16'hB205] = 8'hA9;
mem[16'hB206] = 8'hAA;
mem[16'hB207] = 8'hAB;
mem[16'hB208] = 8'hA4;
mem[16'hB209] = 8'hA5;
mem[16'hB20A] = 8'hA6;
mem[16'hB20B] = 8'hA7;
mem[16'hB20C] = 8'hA0;
mem[16'hB20D] = 8'hA1;
mem[16'hB20E] = 8'hA2;
mem[16'hB20F] = 8'hA3;
mem[16'hB210] = 8'h9C;
mem[16'hB211] = 8'hDD;
mem[16'hB212] = 8'hBE;
mem[16'hB213] = 8'hBF;
mem[16'hB214] = 8'hB8;
mem[16'hB215] = 8'hB9;
mem[16'hB216] = 8'hBA;
mem[16'hB217] = 8'hBB;
mem[16'hB218] = 8'hB4;
mem[16'hB219] = 8'hB5;
mem[16'hB21A] = 8'hB6;
mem[16'hB21B] = 8'hB7;
mem[16'hB21C] = 8'hB0;
mem[16'hB21D] = 8'hB1;
mem[16'hB21E] = 8'hB2;
mem[16'hB21F] = 8'hB3;
mem[16'hB220] = 8'h88;
mem[16'hB221] = 8'h81;
mem[16'hB222] = 8'h8E;
mem[16'hB223] = 8'h8F;
mem[16'hB224] = 8'h88;
mem[16'hB225] = 8'h89;
mem[16'hB226] = 8'h8A;
mem[16'hB227] = 8'h8B;
mem[16'hB228] = 8'h84;
mem[16'hB229] = 8'h85;
mem[16'hB22A] = 8'h86;
mem[16'hB22B] = 8'h87;
mem[16'hB22C] = 8'h80;
mem[16'hB22D] = 8'h81;
mem[16'hB22E] = 8'h82;
mem[16'hB22F] = 8'h83;
mem[16'hB230] = 8'h9C;
mem[16'hB231] = 8'h9D;
mem[16'hB232] = 8'h9E;
mem[16'hB233] = 8'h9F;
mem[16'hB234] = 8'h98;
mem[16'hB235] = 8'h99;
mem[16'hB236] = 8'h9A;
mem[16'hB237] = 8'h9B;
mem[16'hB238] = 8'h94;
mem[16'hB239] = 8'h95;
mem[16'hB23A] = 8'h96;
mem[16'hB23B] = 8'h97;
mem[16'hB23C] = 8'h90;
mem[16'hB23D] = 8'h91;
mem[16'hB23E] = 8'h92;
mem[16'hB23F] = 8'h93;
mem[16'hB240] = 8'hCC;
mem[16'hB241] = 8'h8D;
mem[16'hB242] = 8'hEE;
mem[16'hB243] = 8'hEF;
mem[16'hB244] = 8'hE8;
mem[16'hB245] = 8'hE9;
mem[16'hB246] = 8'hEA;
mem[16'hB247] = 8'hEB;
mem[16'hB248] = 8'hE4;
mem[16'hB249] = 8'hE5;
mem[16'hB24A] = 8'hE6;
mem[16'hB24B] = 8'hE7;
mem[16'hB24C] = 8'hE0;
mem[16'hB24D] = 8'hE1;
mem[16'hB24E] = 8'hE2;
mem[16'hB24F] = 8'hE3;
mem[16'hB250] = 8'hFC;
mem[16'hB251] = 8'hFD;
mem[16'hB252] = 8'hFE;
mem[16'hB253] = 8'hFF;
mem[16'hB254] = 8'hF8;
mem[16'hB255] = 8'hF9;
mem[16'hB256] = 8'hFA;
mem[16'hB257] = 8'hFB;
mem[16'hB258] = 8'hF4;
mem[16'hB259] = 8'hF5;
mem[16'hB25A] = 8'hF6;
mem[16'hB25B] = 8'hF7;
mem[16'hB25C] = 8'hF0;
mem[16'hB25D] = 8'hF1;
mem[16'hB25E] = 8'hF2;
mem[16'hB25F] = 8'hF3;
mem[16'hB260] = 8'hCC;
mem[16'hB261] = 8'hCD;
mem[16'hB262] = 8'hCE;
mem[16'hB263] = 8'hCF;
mem[16'hB264] = 8'hC8;
mem[16'hB265] = 8'hC9;
mem[16'hB266] = 8'hCA;
mem[16'hB267] = 8'hCB;
mem[16'hB268] = 8'hC4;
mem[16'hB269] = 8'hC5;
mem[16'hB26A] = 8'hC6;
mem[16'hB26B] = 8'hC7;
mem[16'hB26C] = 8'hC0;
mem[16'hB26D] = 8'hC1;
mem[16'hB26E] = 8'hC2;
mem[16'hB26F] = 8'hC3;
mem[16'hB270] = 8'hDC;
mem[16'hB271] = 8'hDD;
mem[16'hB272] = 8'hDE;
mem[16'hB273] = 8'hDF;
mem[16'hB274] = 8'hD8;
mem[16'hB275] = 8'hD9;
mem[16'hB276] = 8'hDA;
mem[16'hB277] = 8'hDB;
mem[16'hB278] = 8'hD4;
mem[16'hB279] = 8'hD5;
mem[16'hB27A] = 8'hD6;
mem[16'hB27B] = 8'hD7;
mem[16'hB27C] = 8'hD0;
mem[16'hB27D] = 8'hD1;
mem[16'hB27E] = 8'hD2;
mem[16'hB27F] = 8'hD3;
mem[16'hB280] = 8'h2C;
mem[16'hB281] = 8'h2D;
mem[16'hB282] = 8'h2E;
mem[16'hB283] = 8'h2F;
mem[16'hB284] = 8'h28;
mem[16'hB285] = 8'h29;
mem[16'hB286] = 8'h2A;
mem[16'hB287] = 8'h2B;
mem[16'hB288] = 8'h24;
mem[16'hB289] = 8'h25;
mem[16'hB28A] = 8'h26;
mem[16'hB28B] = 8'h27;
mem[16'hB28C] = 8'h20;
mem[16'hB28D] = 8'h21;
mem[16'hB28E] = 8'h22;
mem[16'hB28F] = 8'h23;
mem[16'hB290] = 8'h3C;
mem[16'hB291] = 8'h3D;
mem[16'hB292] = 8'h3E;
mem[16'hB293] = 8'h3F;
mem[16'hB294] = 8'h38;
mem[16'hB295] = 8'h39;
mem[16'hB296] = 8'h3A;
mem[16'hB297] = 8'h3B;
mem[16'hB298] = 8'h34;
mem[16'hB299] = 8'h35;
mem[16'hB29A] = 8'h36;
mem[16'hB29B] = 8'h37;
mem[16'hB29C] = 8'h30;
mem[16'hB29D] = 8'h31;
mem[16'hB29E] = 8'h32;
mem[16'hB29F] = 8'h33;
mem[16'hB2A0] = 8'h0C;
mem[16'hB2A1] = 8'h0D;
mem[16'hB2A2] = 8'h0E;
mem[16'hB2A3] = 8'h0F;
mem[16'hB2A4] = 8'h08;
mem[16'hB2A5] = 8'h09;
mem[16'hB2A6] = 8'h0A;
mem[16'hB2A7] = 8'h0B;
mem[16'hB2A8] = 8'h04;
mem[16'hB2A9] = 8'h05;
mem[16'hB2AA] = 8'h06;
mem[16'hB2AB] = 8'h07;
mem[16'hB2AC] = 8'h00;
mem[16'hB2AD] = 8'h01;
mem[16'hB2AE] = 8'h02;
mem[16'hB2AF] = 8'h03;
mem[16'hB2B0] = 8'h1C;
mem[16'hB2B1] = 8'h1D;
mem[16'hB2B2] = 8'h1E;
mem[16'hB2B3] = 8'h1F;
mem[16'hB2B4] = 8'h18;
mem[16'hB2B5] = 8'h19;
mem[16'hB2B6] = 8'h1A;
mem[16'hB2B7] = 8'h1B;
mem[16'hB2B8] = 8'h14;
mem[16'hB2B9] = 8'h15;
mem[16'hB2BA] = 8'h16;
mem[16'hB2BB] = 8'h17;
mem[16'hB2BC] = 8'h10;
mem[16'hB2BD] = 8'h11;
mem[16'hB2BE] = 8'h12;
mem[16'hB2BF] = 8'h13;
mem[16'hB2C0] = 8'h6C;
mem[16'hB2C1] = 8'h6D;
mem[16'hB2C2] = 8'h6E;
mem[16'hB2C3] = 8'h6F;
mem[16'hB2C4] = 8'h68;
mem[16'hB2C5] = 8'h69;
mem[16'hB2C6] = 8'h6A;
mem[16'hB2C7] = 8'h6B;
mem[16'hB2C8] = 8'h64;
mem[16'hB2C9] = 8'h65;
mem[16'hB2CA] = 8'h66;
mem[16'hB2CB] = 8'h67;
mem[16'hB2CC] = 8'h60;
mem[16'hB2CD] = 8'h61;
mem[16'hB2CE] = 8'h62;
mem[16'hB2CF] = 8'h63;
mem[16'hB2D0] = 8'h7C;
mem[16'hB2D1] = 8'h7D;
mem[16'hB2D2] = 8'h7E;
mem[16'hB2D3] = 8'h7F;
mem[16'hB2D4] = 8'h78;
mem[16'hB2D5] = 8'h79;
mem[16'hB2D6] = 8'h7A;
mem[16'hB2D7] = 8'h7B;
mem[16'hB2D8] = 8'h74;
mem[16'hB2D9] = 8'h75;
mem[16'hB2DA] = 8'h76;
mem[16'hB2DB] = 8'h77;
mem[16'hB2DC] = 8'h70;
mem[16'hB2DD] = 8'h71;
mem[16'hB2DE] = 8'h72;
mem[16'hB2DF] = 8'h73;
mem[16'hB2E0] = 8'hEC;
mem[16'hB2E1] = 8'h42;
mem[16'hB2E2] = 8'hF7;
mem[16'hB2E3] = 8'h5F;
mem[16'hB2E4] = 8'hE8;
mem[16'hB2E5] = 8'hD0;
mem[16'hB2E6] = 8'hAA;
mem[16'hB2E7] = 8'hFF;
mem[16'hB2E8] = 8'hED;
mem[16'hB2E9] = 8'hBA;
mem[16'hB2EA] = 8'hDF;
mem[16'hB2EB] = 8'hB7;
mem[16'hB2EC] = 8'hF4;
mem[16'hB2ED] = 8'hC9;
mem[16'hB2EE] = 8'h52;
mem[16'hB2EF] = 8'hB1;
mem[16'hB2F0] = 8'hF9;
mem[16'hB2F1] = 8'h57;
mem[16'hB2F2] = 8'h14;
mem[16'hB2F3] = 8'h15;
mem[16'hB2F4] = 8'h12;
mem[16'hB2F5] = 8'hF3;
mem[16'hB2F6] = 8'hF3;
mem[16'hB2F7] = 8'h5B;
mem[16'hB2F8] = 8'hC9;
mem[16'hB2F9] = 8'hA5;
mem[16'hB2FA] = 8'hE2;
mem[16'hB2FB] = 8'hD2;
mem[16'hB2FC] = 8'hAF;
mem[16'hB2FD] = 8'hF7;
mem[16'hB2FE] = 8'hAD;
mem[16'hB2FF] = 8'hFE;
mem[16'hB300] = 8'h5C;
mem[16'hB301] = 8'h1E;
mem[16'hB302] = 8'h2B;
mem[16'hB303] = 8'hBB;
mem[16'hB304] = 8'h05;
mem[16'hB305] = 8'h58;
mem[16'hB306] = 8'h19;
mem[16'hB307] = 8'h2E;
mem[16'hB308] = 8'hB1;
mem[16'hB309] = 8'hE3;
mem[16'hB30A] = 8'hB3;
mem[16'hB30B] = 8'hC1;
mem[16'hB30C] = 8'hB4;
mem[16'hB30D] = 8'h6B;
mem[16'hB30E] = 8'hB2;
mem[16'hB30F] = 8'h5A;
mem[16'hB310] = 8'h2C;
mem[16'hB311] = 8'hF8;
mem[16'hB312] = 8'h18;
mem[16'hB313] = 8'h40;
mem[16'hB314] = 8'h05;
mem[16'hB315] = 8'h79;
mem[16'hB316] = 8'h09;
mem[16'hB317] = 8'hF3;
mem[16'hB318] = 8'h79;
mem[16'hB319] = 8'hE2;
mem[16'hB31A] = 8'h76;
mem[16'hB31B] = 8'hBD;
mem[16'hB31C] = 8'h20;
mem[16'hB31D] = 8'hB2;
mem[16'hB31E] = 8'h7F;
mem[16'hB31F] = 8'hE5;
mem[16'hB320] = 8'h4C;
mem[16'hB321] = 8'h40;
mem[16'hB322] = 8'hDD;
mem[16'hB323] = 8'h4F;
mem[16'hB324] = 8'h82;
mem[16'hB325] = 8'h19;
mem[16'hB326] = 8'h89;
mem[16'hB327] = 8'h46;
mem[16'hB328] = 8'hD6;
mem[16'hB329] = 8'h45;
mem[16'hB32A] = 8'h4B;
mem[16'hB32B] = 8'hD3;
mem[16'hB32C] = 8'h40;
mem[16'hB32D] = 8'h8B;
mem[16'hB32E] = 8'h12;
mem[16'hB32F] = 8'h80;
mem[16'hB330] = 8'h51;
mem[16'hB331] = 8'hC8;
mem[16'hB332] = 8'h5E;
mem[16'hB333] = 8'h52;
mem[16'hB334] = 8'hC8;
mem[16'hB335] = 8'h59;
mem[16'hB336] = 8'h90;
mem[16'hB337] = 8'h0B;
mem[16'hB338] = 8'h97;
mem[16'hB339] = 8'h58;
mem[16'hB33A] = 8'hC7;
mem[16'hB33B] = 8'h57;
mem[16'hB33C] = 8'hF8;
mem[16'hB33D] = 8'hB8;
mem[16'hB33E] = 8'h9D;
mem[16'hB33F] = 8'h1E;
mem[16'hB340] = 8'hEA;
mem[16'hB341] = 8'h4D;
mem[16'hB342] = 8'h47;
mem[16'hB343] = 8'hEE;
mem[16'hB344] = 8'h65;
mem[16'hB345] = 8'hEB;
mem[16'hB346] = 8'h4A;
mem[16'hB347] = 8'h42;
mem[16'hB348] = 8'hE1;
mem[16'hB349] = 8'h68;
mem[16'hB34A] = 8'hE1;
mem[16'hB34B] = 8'h47;
mem[16'hB34C] = 8'hC0;
mem[16'hB34D] = 8'hE1;
mem[16'hB34E] = 8'h59;
mem[16'hB34F] = 8'h4E;
mem[16'hB350] = 8'hF4;
mem[16'hB351] = 8'h5D;
mem[16'hB352] = 8'h0E;
mem[16'hB353] = 8'hFC;
mem[16'hB354] = 8'hB4;
mem[16'hB355] = 8'h5B;
mem[16'hB356] = 8'h42;
mem[16'hB357] = 8'h1D;
mem[16'hB358] = 8'h0B;
mem[16'hB359] = 8'h50;
mem[16'hB35A] = 8'h09;
mem[16'hB35B] = 8'h3E;
mem[16'hB35C] = 8'hE0;
mem[16'hB35D] = 8'h61;
mem[16'hB35E] = 8'h6C;
mem[16'hB35F] = 8'h5E;
mem[16'hB360] = 8'h1C;
mem[16'hB361] = 8'h7E;
mem[16'hB362] = 8'h4B;
mem[16'hB363] = 8'hDF;
mem[16'hB364] = 8'h65;
mem[16'hB365] = 8'h18;
mem[16'hB366] = 8'h79;
mem[16'hB367] = 8'h4E;
mem[16'hB368] = 8'hD5;
mem[16'hB369] = 8'h6C;
mem[16'hB36A] = 8'hD6;
mem[16'hB36B] = 8'h42;
mem[16'hB36C] = 8'hD4;
mem[16'hB36D] = 8'h68;
mem[16'hB36E] = 8'h2E;
mem[16'hB36F] = 8'h46;
mem[16'hB370] = 8'hC9;
mem[16'hB371] = 8'h74;
mem[16'hB372] = 8'h27;
mem[16'hB373] = 8'h5A;
mem[16'hB374] = 8'hCE;
mem[16'hB375] = 8'h70;
mem[16'hB376] = 8'h6E;
mem[16'hB377] = 8'h93;
mem[16'hB378] = 8'h7D;
mem[16'hB379] = 8'h68;
mem[16'hB37A] = 8'h9E;
mem[16'hB37B] = 8'h9B;
mem[16'hB37C] = 8'hAA;
mem[16'hB37D] = 8'h65;
mem[16'hB37E] = 8'hD2;
mem[16'hB37F] = 8'hD3;
mem[16'hB380] = 8'h2D;
mem[16'hB381] = 8'h2D;
mem[16'hB382] = 8'h2E;
mem[16'hB383] = 8'h2F;
mem[16'hB384] = 8'h28;
mem[16'hB385] = 8'h29;
mem[16'hB386] = 8'h2A;
mem[16'hB387] = 8'h2B;
mem[16'hB388] = 8'h24;
mem[16'hB389] = 8'h25;
mem[16'hB38A] = 8'h26;
mem[16'hB38B] = 8'h27;
mem[16'hB38C] = 8'h20;
mem[16'hB38D] = 8'h21;
mem[16'hB38E] = 8'h22;
mem[16'hB38F] = 8'h23;
mem[16'hB390] = 8'h38;
mem[16'hB391] = 8'h3D;
mem[16'hB392] = 8'h3E;
mem[16'hB393] = 8'h3F;
mem[16'hB394] = 8'h38;
mem[16'hB395] = 8'h39;
mem[16'hB396] = 8'h3A;
mem[16'hB397] = 8'h3B;
mem[16'hB398] = 8'h34;
mem[16'hB399] = 8'h35;
mem[16'hB39A] = 8'h36;
mem[16'hB39B] = 8'h37;
mem[16'hB39C] = 8'h30;
mem[16'hB39D] = 8'h31;
mem[16'hB39E] = 8'h32;
mem[16'hB39F] = 8'h33;
mem[16'hB3A0] = 8'h2F;
mem[16'hB3A1] = 8'h0D;
mem[16'hB3A2] = 8'h0E;
mem[16'hB3A3] = 8'h0F;
mem[16'hB3A4] = 8'h08;
mem[16'hB3A5] = 8'h09;
mem[16'hB3A6] = 8'h0A;
mem[16'hB3A7] = 8'h0B;
mem[16'hB3A8] = 8'h04;
mem[16'hB3A9] = 8'h05;
mem[16'hB3AA] = 8'h06;
mem[16'hB3AB] = 8'h07;
mem[16'hB3AC] = 8'h00;
mem[16'hB3AD] = 8'h01;
mem[16'hB3AE] = 8'h02;
mem[16'hB3AF] = 8'h03;
mem[16'hB3B0] = 8'h1D;
mem[16'hB3B1] = 8'h1D;
mem[16'hB3B2] = 8'h1E;
mem[16'hB3B3] = 8'h1F;
mem[16'hB3B4] = 8'h18;
mem[16'hB3B5] = 8'h19;
mem[16'hB3B6] = 8'h1A;
mem[16'hB3B7] = 8'h1B;
mem[16'hB3B8] = 8'h14;
mem[16'hB3B9] = 8'h15;
mem[16'hB3BA] = 8'h16;
mem[16'hB3BB] = 8'h17;
mem[16'hB3BC] = 8'h10;
mem[16'hB3BD] = 8'h11;
mem[16'hB3BE] = 8'h12;
mem[16'hB3BF] = 8'h13;
mem[16'hB3C0] = 8'hFD;
mem[16'hB3C1] = 8'h6D;
mem[16'hB3C2] = 8'h6E;
mem[16'hB3C3] = 8'h6F;
mem[16'hB3C4] = 8'h68;
mem[16'hB3C5] = 8'h69;
mem[16'hB3C6] = 8'h6A;
mem[16'hB3C7] = 8'h6B;
mem[16'hB3C8] = 8'h64;
mem[16'hB3C9] = 8'h65;
mem[16'hB3CA] = 8'h66;
mem[16'hB3CB] = 8'h67;
mem[16'hB3CC] = 8'h60;
mem[16'hB3CD] = 8'h61;
mem[16'hB3CE] = 8'h62;
mem[16'hB3CF] = 8'h63;
mem[16'hB3D0] = 8'h7C;
mem[16'hB3D1] = 8'hE1;
mem[16'hB3D2] = 8'hD6;
mem[16'hB3D3] = 8'h7F;
mem[16'hB3D4] = 8'hD8;
mem[16'hB3D5] = 8'h79;
mem[16'hB3D6] = 8'h7A;
mem[16'hB3D7] = 8'h7B;
mem[16'hB3D8] = 8'h74;
mem[16'hB3D9] = 8'h75;
mem[16'hB3DA] = 8'h76;
mem[16'hB3DB] = 8'h77;
mem[16'hB3DC] = 8'h70;
mem[16'hB3DD] = 8'h71;
mem[16'hB3DE] = 8'h72;
mem[16'hB3DF] = 8'h73;
mem[16'hB3E0] = 8'h4C;
mem[16'hB3E1] = 8'h4D;
mem[16'hB3E2] = 8'h4E;
mem[16'hB3E3] = 8'h4F;
mem[16'hB3E4] = 8'h48;
mem[16'hB3E5] = 8'h49;
mem[16'hB3E6] = 8'h4A;
mem[16'hB3E7] = 8'h4B;
mem[16'hB3E8] = 8'h44;
mem[16'hB3E9] = 8'h45;
mem[16'hB3EA] = 8'h46;
mem[16'hB3EB] = 8'h47;
mem[16'hB3EC] = 8'h40;
mem[16'hB3ED] = 8'h41;
mem[16'hB3EE] = 8'h42;
mem[16'hB3EF] = 8'h43;
mem[16'hB3F0] = 8'h5D;
mem[16'hB3F1] = 8'h5D;
mem[16'hB3F2] = 8'h5F;
mem[16'hB3F3] = 8'h5C;
mem[16'hB3F4] = 8'h59;
mem[16'hB3F5] = 8'h59;
mem[16'hB3F6] = 8'h5A;
mem[16'hB3F7] = 8'h5B;
mem[16'hB3F8] = 8'h54;
mem[16'hB3F9] = 8'h55;
mem[16'hB3FA] = 8'h56;
mem[16'hB3FB] = 8'h57;
mem[16'hB3FC] = 8'h50;
mem[16'hB3FD] = 8'h51;
mem[16'hB3FE] = 8'h52;
mem[16'hB3FF] = 8'h53;
mem[16'hB400] = 8'h08;
mem[16'hB401] = 8'h30;
mem[16'hB402] = 8'h01;
mem[16'hB403] = 8'h4C;
mem[16'hB404] = 8'hD0;
mem[16'hB405] = 8'h01;
mem[16'hB406] = 8'h4C;
mem[16'hB407] = 8'h8A;
mem[16'hB408] = 8'h48;
mem[16'hB409] = 8'h98;
mem[16'hB40A] = 8'h48;
mem[16'hB40B] = 8'hA2;
mem[16'hB40C] = 8'h1F;
mem[16'hB40D] = 8'hB5;
mem[16'hB40E] = 8'h00;
mem[16'hB40F] = 8'h9D;
mem[16'hB410] = 8'hC0;
mem[16'hB411] = 8'hB4;
mem[16'hB412] = 8'hCA;
mem[16'hB413] = 8'h10;
mem[16'hB414] = 8'hF8;
mem[16'hB415] = 8'h20;
mem[16'hB416] = 8'h68;
mem[16'hB417] = 8'hB4;
mem[16'hB418] = 8'hAD;
mem[16'hB419] = 8'h07;
mem[16'hB41A] = 8'hA0;
mem[16'hB41B] = 8'h20;
mem[16'hB41C] = 8'h00;
mem[16'hB41D] = 8'hBB;
mem[16'hB41E] = 8'h20;
mem[16'hB41F] = 8'h68;
mem[16'hB420] = 8'hB4;
mem[16'hB421] = 8'hA2;
mem[16'hB422] = 8'h1F;
mem[16'hB423] = 8'hBD;
mem[16'hB424] = 8'hC0;
mem[16'hB425] = 8'hB4;
mem[16'hB426] = 8'h95;
mem[16'hB427] = 8'h00;
mem[16'hB428] = 8'hCA;
mem[16'hB429] = 8'h10;
mem[16'hB42A] = 8'hF8;
mem[16'hB42B] = 8'hA9;
mem[16'hB42C] = 8'h85;
mem[16'hB42D] = 8'h8D;
mem[16'hB42E] = 8'h00;
mem[16'hB42F] = 8'hA8;
mem[16'hB430] = 8'hA9;
mem[16'hB431] = 8'hA9;
mem[16'hB432] = 8'h8D;
mem[16'hB433] = 8'h01;
mem[16'hB434] = 8'hA8;
mem[16'hB435] = 8'hA9;
mem[16'hB436] = 8'hB3;
mem[16'hB437] = 8'h8D;
mem[16'hB438] = 8'h02;
mem[16'hB439] = 8'hA8;
mem[16'hB43A] = 8'hAD;
mem[16'hB43B] = 8'h08;
mem[16'hB43C] = 8'hB4;
mem[16'hB43D] = 8'h8D;
mem[16'hB43E] = 8'h03;
mem[16'hB43F] = 8'hA8;
mem[16'hB440] = 8'hA9;
mem[16'hB441] = 8'hA9;
mem[16'hB442] = 8'h8D;
mem[16'hB443] = 8'h04;
mem[16'hB444] = 8'hA8;
mem[16'hB445] = 8'hA9;
mem[16'hB446] = 8'hFF;
mem[16'hB447] = 8'h8D;
mem[16'hB448] = 8'h05;
mem[16'hB449] = 8'hA8;
mem[16'hB44A] = 8'hAD;
mem[16'hB44B] = 8'h08;
mem[16'hB44C] = 8'hB4;
mem[16'hB44D] = 8'h8D;
mem[16'hB44E] = 8'h06;
mem[16'hB44F] = 8'hA8;
mem[16'hB450] = 8'hA9;
mem[16'hB451] = 8'h60;
mem[16'hB452] = 8'h8D;
mem[16'hB453] = 8'h07;
mem[16'hB454] = 8'hA8;
mem[16'hB455] = 8'h68;
mem[16'hB456] = 8'hA8;
mem[16'hB457] = 8'h68;
mem[16'hB458] = 8'hAA;
mem[16'hB459] = 8'hAD;
mem[16'hB45A] = 8'h08;
mem[16'hB45B] = 8'hA0;
mem[16'hB45C] = 8'hC9;
mem[16'hB45D] = 8'h01;
mem[16'hB45E] = 8'h90;
mem[16'hB45F] = 8'h04;
mem[16'hB460] = 8'h28;
mem[16'hB461] = 8'h38;
mem[16'hB462] = 8'h60;
mem[16'hB463] = 8'h20;
mem[16'hB464] = 8'h28;
mem[16'hB465] = 8'h18;
mem[16'hB466] = 8'h60;
mem[16'hB467] = 8'h20;
mem[16'hB468] = 8'hAE;
mem[16'hB469] = 8'h07;
mem[16'hB46A] = 8'hA0;
mem[16'hB46B] = 8'hBD;
mem[16'hB46C] = 8'hA0;
mem[16'hB46D] = 8'hB4;
mem[16'hB46E] = 8'h85;
mem[16'hB46F] = 8'h14;
mem[16'hB470] = 8'hBD;
mem[16'hB471] = 8'hAA;
mem[16'hB472] = 8'hB4;
mem[16'hB473] = 8'h85;
mem[16'hB474] = 8'h15;
mem[16'hB475] = 8'hBD;
mem[16'hB476] = 8'hB4;
mem[16'hB477] = 8'hB4;
mem[16'hB478] = 8'h85;
mem[16'hB479] = 8'h16;
mem[16'hB47A] = 8'hA0;
mem[16'hB47B] = 8'h00;
mem[16'hB47C] = 8'h84;
mem[16'hB47D] = 8'h08;
mem[16'hB47E] = 8'hA9;
mem[16'hB47F] = 8'hA8;
mem[16'hB480] = 8'h85;
mem[16'hB481] = 8'h09;
mem[16'hB482] = 8'h46;
mem[16'hB483] = 8'h16;
mem[16'hB484] = 8'h66;
mem[16'hB485] = 8'h15;
mem[16'hB486] = 8'h66;
mem[16'hB487] = 8'h14;
mem[16'hB488] = 8'h90;
mem[16'hB489] = 8'h0D;
mem[16'hB48A] = 8'hB0;
mem[16'hB48B] = 8'h01;
mem[16'hB48C] = 8'h4C;
mem[16'hB48D] = 8'h98;
mem[16'hB48E] = 8'h49;
mem[16'hB48F] = 8'hAC;
mem[16'hB490] = 8'h51;
mem[16'hB491] = 8'h08;
mem[16'hB492] = 8'h91;
mem[16'hB493] = 8'h08;
mem[16'hB494] = 8'hC8;
mem[16'hB495] = 8'hD0;
mem[16'hB496] = 8'hF6;
mem[16'hB497] = 8'hE6;
mem[16'hB498] = 8'h09;
mem[16'hB499] = 8'hA5;
mem[16'hB49A] = 8'h09;
mem[16'hB49B] = 8'hC9;
mem[16'hB49C] = 8'hC0;
mem[16'hB49D] = 8'hD0;
mem[16'hB49E] = 8'hE3;
mem[16'hB49F] = 8'h60;
mem[16'hB4A0] = 8'h00;
mem[16'hB4A1] = 8'h10;
mem[16'hB4A2] = 8'h10;
mem[16'hB4A3] = 8'h10;
mem[16'hB4A4] = 8'h10;
mem[16'hB4A5] = 8'h10;
mem[16'hB4A6] = 8'h10;
mem[16'hB4A7] = 8'h10;
mem[16'hB4A8] = 8'h00;
mem[16'hB4A9] = 8'h00;
mem[16'hB4AA] = 8'h60;
mem[16'hB4AB] = 8'hE0;
mem[16'hB4AC] = 8'h60;
mem[16'hB4AD] = 8'hE0;
mem[16'hB4AE] = 8'h60;
mem[16'hB4AF] = 8'hEC;
mem[16'hB4B0] = 8'h6C;
mem[16'hB4B1] = 8'hEC;
mem[16'hB4B2] = 8'h00;
mem[16'hB4B3] = 8'h00;
mem[16'hB4B4] = 8'hF8;
mem[16'hB4B5] = 8'hF9;
mem[16'hB4B6] = 8'hFF;
mem[16'hB4B7] = 8'hF9;
mem[16'hB4B8] = 8'hFF;
mem[16'hB4B9] = 8'hF9;
mem[16'hB4BA] = 8'hFF;
mem[16'hB4BB] = 8'hF9;
mem[16'hB4BC] = 8'hF8;
mem[16'hB4BD] = 8'hF8;
mem[16'hB4BE] = 8'hA9;
mem[16'hB4BF] = 8'h08;
mem[16'hB4C0] = 8'h00;
mem[16'hB4C1] = 8'h9C;
mem[16'hB4C2] = 8'h00;
mem[16'hB4C3] = 8'h08;
mem[16'hB4C4] = 8'h3A;
mem[16'hB4C5] = 8'h03;
mem[16'hB4C6] = 8'h00;
mem[16'hB4C7] = 8'h00;
mem[16'hB4C8] = 8'h00;
mem[16'hB4C9] = 8'hC0;
mem[16'hB4CA] = 8'h60;
mem[16'hB4CB] = 8'h01;
mem[16'hB4CC] = 8'h05;
mem[16'hB4CD] = 8'h00;
mem[16'hB4CE] = 8'h00;
mem[16'hB4CF] = 8'h6B;
mem[16'hB4D0] = 8'h00;
mem[16'hB4D1] = 8'h9C;
mem[16'hB4D2] = 8'h00;
mem[16'hB4D3] = 8'h04;
mem[16'hB4D4] = 8'h00;
mem[16'hB4D5] = 8'h00;
mem[16'hB4D6] = 8'h00;
mem[16'hB4D7] = 8'h00;
mem[16'hB4D8] = 8'hFF;
mem[16'hB4D9] = 8'h0C;
mem[16'hB4DA] = 8'h00;
mem[16'hB4DB] = 8'h56;
mem[16'hB4DC] = 8'hFF;
mem[16'hB4DD] = 8'hFF;
mem[16'hB4DE] = 8'h00;
mem[16'hB4DF] = 8'h00;
mem[16'hB4E0] = 8'h41;
mem[16'hB4E1] = 8'h00;
mem[16'hB4E2] = 8'h00;
mem[16'hB4E3] = 8'h00;
mem[16'hB4E4] = 8'h00;
mem[16'hB4E5] = 8'h00;
mem[16'hB4E6] = 8'hBE;
mem[16'hB4E7] = 8'h00;
mem[16'hB4E8] = 8'h4C;
mem[16'hB4E9] = 8'hC0;
mem[16'hB4EA] = 8'h60;
mem[16'hB4EB] = 8'h00;
mem[16'hB4EC] = 8'hFF;
mem[16'hB4ED] = 8'hAA;
mem[16'hB4EE] = 8'hAC;
mem[16'hB4EF] = 8'h5F;
mem[16'hB4F0] = 8'hFF;
mem[16'hB4F1] = 8'hFF;
mem[16'hB4F2] = 8'hFF;
mem[16'hB4F3] = 8'hFF;
mem[16'hB4F4] = 8'hFF;
mem[16'hB4F5] = 8'hFF;
mem[16'hB4F6] = 8'hFF;
mem[16'hB4F7] = 8'hFF;
mem[16'hB4F8] = 8'hFF;
mem[16'hB4F9] = 8'hFF;
mem[16'hB4FA] = 8'hFF;
mem[16'hB4FB] = 8'hFF;
mem[16'hB4FC] = 8'h0B;
mem[16'hB4FD] = 8'hFF;
mem[16'hB4FE] = 8'hFF;
mem[16'hB4FF] = 8'hFF;
mem[16'hB500] = 8'hE0;
mem[16'hB501] = 8'h40;
mem[16'hB502] = 8'h1B;
mem[16'hB503] = 8'hE3;
mem[16'hB504] = 8'hEB;
mem[16'hB505] = 8'h1F;
mem[16'hB506] = 8'hE6;
mem[16'hB507] = 8'h08;
mem[16'hB508] = 8'h11;
mem[16'hB509] = 8'hE9;
mem[16'hB50A] = 8'hDF;
mem[16'hB50B] = 8'h11;
mem[16'hB50C] = 8'hEC;
mem[16'hB50D] = 8'hF5;
mem[16'hB50E] = 8'h14;
mem[16'hB50F] = 8'h06;
mem[16'hB510] = 8'hBC;
mem[16'hB511] = 8'h94;
mem[16'hB512] = 8'hB9;
mem[16'hB513] = 8'h17;
mem[16'hB514] = 8'hB1;
mem[16'hB515] = 8'hB8;
mem[16'hB516] = 8'hBF;
mem[16'hB517] = 8'hB1;
mem[16'hB518] = 8'h1E;
mem[16'hB519] = 8'h68;
mem[16'hB51A] = 8'h36;
mem[16'hB51B] = 8'h77;
mem[16'hB51C] = 8'h78;
mem[16'hB51D] = 8'h29;
mem[16'hB51E] = 8'hB7;
mem[16'hB51F] = 8'hB9;
mem[16'hB520] = 8'hA5;
mem[16'hB521] = 8'h7A;
mem[16'hB522] = 8'h87;
mem[16'hB523] = 8'h8E;
mem[16'hB524] = 8'h22;
mem[16'hB525] = 8'h34;
mem[16'hB526] = 8'h0A;
mem[16'hB527] = 8'h4B;
mem[16'hB528] = 8'h22;
mem[16'hB529] = 8'h8F;
mem[16'hB52A] = 8'h23;
mem[16'hB52B] = 8'h86;
mem[16'hB52C] = 8'h45;
mem[16'hB52D] = 8'h81;
mem[16'hB52E] = 8'h12;
mem[16'hB52F] = 8'h8D;
mem[16'hB530] = 8'h6C;
mem[16'hB531] = 8'h85;
mem[16'hB532] = 8'hBE;
mem[16'hB533] = 8'hFC;
mem[16'hB534] = 8'h2D;
mem[16'hB535] = 8'h30;
mem[16'hB536] = 8'h89;
mem[16'hB537] = 8'hBB;
mem[16'hB538] = 8'h10;
mem[16'hB539] = 8'h20;
mem[16'hB53A] = 8'hDA;
mem[16'hB53B] = 8'hBD;
mem[16'hB53C] = 8'h25;
mem[16'hB53D] = 8'h54;
mem[16'hB53E] = 8'hB2;
mem[16'hB53F] = 8'hE3;
mem[16'hB540] = 8'h59;
mem[16'hB541] = 8'h44;
mem[16'hB542] = 8'hFD;
mem[16'hB543] = 8'hCF;
mem[16'hB544] = 8'h6C;
mem[16'hB545] = 8'h5C;
mem[16'hB546] = 8'hA6;
mem[16'hB547] = 8'hC1;
mem[16'hB548] = 8'h51;
mem[16'hB549] = 8'h80;
mem[16'hB54A] = 8'h43;
mem[16'hB54B] = 8'hE0;
mem[16'hB54C] = 8'hC9;
mem[16'hB54D] = 8'hE3;
mem[16'hB54E] = 8'h12;
mem[16'hB54F] = 8'hF2;
mem[16'hB550] = 8'h55;
mem[16'hB551] = 8'hAD;
mem[16'hB552] = 8'hDE;
mem[16'hB553] = 8'h7B;
mem[16'hB554] = 8'h4D;
mem[16'hB555] = 8'h44;
mem[16'hB556] = 8'h7A;
mem[16'hB557] = 8'h3B;
mem[16'hB558] = 8'h49;
mem[16'hB559] = 8'h77;
mem[16'hB55A] = 8'h36;
mem[16'hB55B] = 8'h4A;
mem[16'hB55C] = 8'h74;
mem[16'hB55D] = 8'h31;
mem[16'hB55E] = 8'h4F;
mem[16'hB55F] = 8'h75;
mem[16'hB560] = 8'h0C;
mem[16'hB561] = 8'hAD;
mem[16'hB562] = 8'h4B;
mem[16'hB563] = 8'h29;
mem[16'hB564] = 8'hC8;
mem[16'hB565] = 8'h6C;
mem[16'hB566] = 8'hCA;
mem[16'hB567] = 8'hE2;
mem[16'hB568] = 8'hC3;
mem[16'hB569] = 8'h6F;
mem[16'hB56A] = 8'h7B;
mem[16'hB56B] = 8'h5C;
mem[16'hB56C] = 8'h75;
mem[16'hB56D] = 8'hD1;
mem[16'hB56E] = 8'hC9;
mem[16'hB56F] = 8'h6A;
mem[16'hB570] = 8'h1A;
mem[16'hB571] = 8'hDD;
mem[16'hB572] = 8'h7B;
mem[16'hB573] = 8'hDF;
mem[16'hB574] = 8'hF1;
mem[16'hB575] = 8'hDE;
mem[16'hB576] = 8'h70;
mem[16'hB577] = 8'h66;
mem[16'hB578] = 8'h47;
mem[16'hB579] = 8'h60;
mem[16'hB57A] = 8'hD3;
mem[16'hB57B] = 8'hDD;
mem[16'hB57C] = 8'h7A;
mem[16'hB57D] = 8'h6C;
mem[16'hB57E] = 8'h52;
mem[16'hB57F] = 8'h13;
mem[16'hB580] = 8'h8A;
mem[16'hB581] = 8'h27;
mem[16'hB582] = 8'h4E;
mem[16'hB583] = 8'hE6;
mem[16'hB584] = 8'hAD;
mem[16'hB585] = 8'h27;
mem[16'hB586] = 8'h83;
mem[16'hB587] = 8'h3E;
mem[16'hB588] = 8'hA1;
mem[16'hB589] = 8'h2D;
mem[16'hB58A] = 8'hE0;
mem[16'hB58B] = 8'h2F;
mem[16'hB58C] = 8'hF0;
mem[16'hB58D] = 8'hDD;
mem[16'hB58E] = 8'hE4;
mem[16'hB58F] = 8'h2D;
mem[16'hB590] = 8'hEC;
mem[16'hB591] = 8'hC9;
mem[16'hB592] = 8'h5E;
mem[16'hB593] = 8'h3D;
mem[16'hB594] = 8'h39;
mem[16'hB595] = 8'h3D;
mem[16'hB596] = 8'h39;
mem[16'hB597] = 8'h3D;
mem[16'hB598] = 8'h31;
mem[16'hB599] = 8'h35;
mem[16'hB59A] = 8'h31;
mem[16'hB59B] = 8'h31;
mem[16'hB59C] = 8'h33;
mem[16'hB59D] = 8'h31;
mem[16'hB59E] = 8'h37;
mem[16'hB59F] = 8'h31;
mem[16'hB5A0] = 8'h0B;
mem[16'hB5A1] = 8'h09;
mem[16'hB5A2] = 8'h0F;
mem[16'hB5A3] = 8'hA6;
mem[16'hB5A4] = 8'h08;
mem[16'hB5A5] = 8'h8C;
mem[16'hB5A6] = 8'h1A;
mem[16'hB5A7] = 8'hA2;
mem[16'hB5A8] = 8'h44;
mem[16'hB5A9] = 8'h80;
mem[16'hB5AA] = 8'h17;
mem[16'hB5AB] = 8'hA2;
mem[16'hB5AC] = 8'h07;
mem[16'hB5AD] = 8'h28;
mem[16'hB5AE] = 8'h07;
mem[16'hB5AF] = 8'hD3;
mem[16'hB5B0] = 8'h14;
mem[16'hB5B1] = 8'hB4;
mem[16'hB5B2] = 8'h3E;
mem[16'hB5B3] = 8'h9A;
mem[16'hB5B4] = 8'h08;
mem[16'hB5B5] = 8'hB0;
mem[16'hB5B6] = 8'h1B;
mem[16'hB5B7] = 8'h9E;
mem[16'hB5B8] = 8'h05;
mem[16'hB5B9] = 8'hB3;
mem[16'hB5BA] = 8'h1C;
mem[16'hB5BB] = 8'hAA;
mem[16'hB5BC] = 8'h9E;
mem[16'hB5BD] = 8'hD1;
mem[16'hB5BE] = 8'hAF;
mem[16'hB5BF] = 8'h9F;
mem[16'hB5C0] = 8'hAC;
mem[16'hB5C1] = 8'h7D;
mem[16'hB5C2] = 8'h95;
mem[16'hB5C3] = 8'hA6;
mem[16'hB5C4] = 8'hFF;
mem[16'hB5C5] = 8'h99;
mem[16'hB5C6] = 8'h7B;
mem[16'hB5C7] = 8'hAD;
mem[16'hB5C8] = 8'h74;
mem[16'hB5C9] = 8'hB5;
mem[16'hB5CA] = 8'h95;
mem[16'hB5CB] = 8'hA1;
mem[16'hB5CC] = 8'h71;
mem[16'hB5CD] = 8'hB1;
mem[16'hB5CE] = 8'h8D;
mem[16'hB5CF] = 8'hCA;
mem[16'hB5D0] = 8'h6D;
mem[16'hB5D1] = 8'hF0;
mem[16'hB5D2] = 8'h76;
mem[16'hB5D3] = 8'hDF;
mem[16'hB5D4] = 8'h10;
mem[16'hB5D5] = 8'h11;
mem[16'hB5D6] = 8'h1A;
mem[16'hB5D7] = 8'hA2;
mem[16'hB5D8] = 8'hD2;
mem[16'hB5D9] = 8'h63;
mem[16'hB5DA] = 8'hCB;
mem[16'hB5DB] = 8'h77;
mem[16'hB5DC] = 8'hDB;
mem[16'hB5DD] = 8'hFC;
mem[16'hB5DE] = 8'h9A;
mem[16'hB5DF] = 8'hC6;
mem[16'hB5E0] = 8'hEA;
mem[16'hB5E1] = 8'h47;
mem[16'hB5E2] = 8'hF3;
mem[16'hB5E3] = 8'hC3;
mem[16'hB5E4] = 8'h88;
mem[16'hB5E5] = 8'h59;
mem[16'hB5E6] = 8'hB1;
mem[16'hB5E7] = 8'h82;
mem[16'hB5E8] = 8'hF6;
mem[16'hB5E9] = 8'h95;
mem[16'hB5EA] = 8'h9E;
mem[16'hB5EB] = 8'h27;
mem[16'hB5EC] = 8'h09;
mem[16'hB5ED] = 8'hE1;
mem[16'hB5EE] = 8'h42;
mem[16'hB5EF] = 8'hC7;
mem[16'hB5F0] = 8'h54;
mem[16'hB5F1] = 8'hF8;
mem[16'hB5F2] = 8'h54;
mem[16'hB5F3] = 8'h15;
mem[16'hB5F4] = 8'h12;
mem[16'hB5F5] = 8'h13;
mem[16'hB5F6] = 8'h10;
mem[16'hB5F7] = 8'h52;
mem[16'hB5F8] = 8'h94;
mem[16'hB5F9] = 8'hD0;
mem[16'hB5FA] = 8'h5F;
mem[16'hB5FB] = 8'hCF;
mem[16'hB5FC] = 8'h01;
mem[16'hB5FD] = 8'h59;
mem[16'hB5FE] = 8'h9A;
mem[16'hB5FF] = 8'h83;
mem[16'hB600] = 8'h57;
mem[16'hB601] = 8'h64;
mem[16'hB602] = 8'h10;
mem[16'hB603] = 8'h5F;
mem[16'hB604] = 8'hAF;
mem[16'hB605] = 8'h00;
mem[16'hB606] = 8'hBF;
mem[16'hB607] = 8'h26;
mem[16'hB608] = 8'hAC;
mem[16'hB609] = 8'h05;
mem[16'hB60A] = 8'hC6;
mem[16'hB60B] = 8'h0E;
mem[16'hB60C] = 8'h06;
mem[16'hB60D] = 8'hAB;
mem[16'hB60E] = 8'h1F;
mem[16'hB60F] = 8'h2A;
mem[16'hB610] = 8'h7C;
mem[16'hB611] = 8'h18;
mem[16'hB612] = 8'hB5;
mem[16'hB613] = 8'h76;
mem[16'hB614] = 8'hB9;
mem[16'hB615] = 8'h69;
mem[16'hB616] = 8'hBD;
mem[16'hB617] = 8'h06;
mem[16'hB618] = 8'h3E;
mem[16'hB619] = 8'h75;
mem[16'hB61A] = 8'hFA;
mem[16'hB61B] = 8'h96;
mem[16'hB61C] = 8'h06;
mem[16'hB61D] = 8'h34;
mem[16'hB61E] = 8'h0F;
mem[16'hB61F] = 8'h38;
mem[16'hB620] = 8'h4C;
mem[16'hB621] = 8'h30;
mem[16'hB622] = 8'h00;
mem[16'hB623] = 8'h4F;
mem[16'hB624] = 8'h35;
mem[16'hB625] = 8'h05;
mem[16'hB626] = 8'h4A;
mem[16'hB627] = 8'h2B;
mem[16'hB628] = 8'h64;
mem[16'hB629] = 8'h4D;
mem[16'hB62A] = 8'h76;
mem[16'hB62B] = 8'h8F;
mem[16'hB62C] = 8'h5D;
mem[16'hB62D] = 8'h0D;
mem[16'hB62E] = 8'h42;
mem[16'hB62F] = 8'h73;
mem[16'hB630] = 8'h64;
mem[16'hB631] = 8'hD1;
mem[16'hB632] = 8'hDF;
mem[16'hB633] = 8'h29;
mem[16'hB634] = 8'h38;
mem[16'hB635] = 8'hF1;
mem[16'hB636] = 8'h33;
mem[16'hB637] = 8'h8F;
mem[16'hB638] = 8'hB4;
mem[16'hB639] = 8'h11;
mem[16'hB63A] = 8'h23;
mem[16'hB63B] = 8'h1F;
mem[16'hB63C] = 8'h40;
mem[16'hB63D] = 8'h69;
mem[16'hB63E] = 8'hB2;
mem[16'hB63F] = 8'h97;
mem[16'hB640] = 8'h57;
mem[16'hB641] = 8'h8D;
mem[16'hB642] = 8'hDF;
mem[16'hB643] = 8'h49;
mem[16'hB644] = 8'hE2;
mem[16'hB645] = 8'h54;
mem[16'hB646] = 8'h64;
mem[16'hB647] = 8'h2B;
mem[16'hB648] = 8'h59;
mem[16'hB649] = 8'h69;
mem[16'hB64A] = 8'h26;
mem[16'hB64B] = 8'h4E;
mem[16'hB64C] = 8'hD0;
mem[16'hB64D] = 8'hC1;
mem[16'hB64E] = 8'h66;
mem[16'hB64F] = 8'h56;
mem[16'hB650] = 8'h41;
mem[16'hB651] = 8'h75;
mem[16'hB652] = 8'h3E;
mem[16'hB653] = 8'h9F;
mem[16'hB654] = 8'h46;
mem[16'hB655] = 8'hF9;
mem[16'hB656] = 8'h56;
mem[16'hB657] = 8'h63;
mem[16'hB658] = 8'h69;
mem[16'hB659] = 8'hF5;
mem[16'hB65A] = 8'h5A;
mem[16'hB65B] = 8'hDE;
mem[16'hB65C] = 8'hFF;
mem[16'hB65D] = 8'h6C;
mem[16'hB65E] = 8'hF2;
mem[16'hB65F] = 8'h5D;
mem[16'hB660] = 8'hE5;
mem[16'hB661] = 8'hCE;
mem[16'hB662] = 8'h53;
mem[16'hB663] = 8'hCF;
mem[16'hB664] = 8'h78;
mem[16'hB665] = 8'h51;
mem[16'hB666] = 8'hC0;
mem[16'hB667] = 8'hC1;
mem[16'hB668] = 8'h59;
mem[16'hB669] = 8'hC5;
mem[16'hB66A] = 8'h77;
mem[16'hB66B] = 8'hEE;
mem[16'hB66C] = 8'h30;
mem[16'hB66D] = 8'h5C;
mem[16'hB66E] = 8'hC2;
mem[16'hB66F] = 8'h6C;
mem[16'hB670] = 8'hF5;
mem[16'hB671] = 8'h1D;
mem[16'hB672] = 8'h43;
mem[16'hB673] = 8'hDF;
mem[16'hB674] = 8'h75;
mem[16'hB675] = 8'h51;
mem[16'hB676] = 8'hCA;
mem[16'hB677] = 8'h07;
mem[16'hB678] = 8'hB4;
mem[16'hB679] = 8'h6B;
mem[16'hB67A] = 8'hD6;
mem[16'hB67B] = 8'h7B;
mem[16'hB67C] = 8'h5A;
mem[16'hB67D] = 8'h48;
mem[16'hB67E] = 8'h92;
mem[16'hB67F] = 8'h7F;
mem[16'hB680] = 8'hB5;
mem[16'hB681] = 8'hAD;
mem[16'hB682] = 8'h82;
mem[16'hB683] = 8'hB6;
mem[16'hB684] = 8'hE8;
mem[16'hB685] = 8'h85;
mem[16'hB686] = 8'hB2;
mem[16'hB687] = 8'h21;
mem[16'hB688] = 8'h2E;
mem[16'hB689] = 8'h0C;
mem[16'hB68A] = 8'hE6;
mem[16'hB68B] = 8'hA2;
mem[16'hB68C] = 8'h30;
mem[16'hB68D] = 8'hB9;
mem[16'hB68E] = 8'h0B;
mem[16'hB68F] = 8'h2C;
mem[16'hB690] = 8'h39;
mem[16'hB691] = 8'h2D;
mem[16'hB692] = 8'hBB;
mem[16'hB693] = 8'h2F;
mem[16'hB694] = 8'hB2;
mem[16'hB695] = 8'h9F;
mem[16'hB696] = 8'h2A;
mem[16'hB697] = 8'hA6;
mem[16'hB698] = 8'h34;
mem[16'hB699] = 8'h9B;
mem[16'hB69A] = 8'h9C;
mem[16'hB69B] = 8'hAF;
mem[16'hB69C] = 8'h3A;
mem[16'hB69D] = 8'h3B;
mem[16'hB69E] = 8'h1B;
mem[16'hB69F] = 8'hC3;
mem[16'hB6A0] = 8'h09;
mem[16'hB6A1] = 8'h1D;
mem[16'hB6A2] = 8'h27;
mem[16'hB6A3] = 8'hFC;
mem[16'hB6A4] = 8'h8D;
mem[16'hB6A5] = 8'h19;
mem[16'hB6A6] = 8'h80;
mem[16'hB6A7] = 8'hAD;
mem[16'hB6A8] = 8'h14;
mem[16'hB6A9] = 8'h98;
mem[16'hB6AA] = 8'h06;
mem[16'hB6AB] = 8'hB7;
mem[16'hB6AC] = 8'hAA;
mem[16'hB6AD] = 8'h99;
mem[16'hB6AE] = 8'h08;
mem[16'hB6AF] = 8'h09;
mem[16'hB6B0] = 8'h99;
mem[16'hB6B1] = 8'h0D;
mem[16'hB6B2] = 8'h94;
mem[16'hB6B3] = 8'hB9;
mem[16'hB6B4] = 8'h08;
mem[16'hB6B5] = 8'h84;
mem[16'hB6B6] = 8'h1A;
mem[16'hB6B7] = 8'hAA;
mem[16'hB6B8] = 8'h89;
mem[16'hB6B9] = 8'h14;
mem[16'hB6BA] = 8'hA7;
mem[16'hB6BB] = 8'h8A;
mem[16'hB6BC] = 8'h12;
mem[16'hB6BD] = 8'hA0;
mem[16'hB6BE] = 8'h8F;
mem[16'hB6BF] = 8'h10;
mem[16'hB6C0] = 8'hDD;
mem[16'hB6C1] = 8'hE5;
mem[16'hB6C2] = 8'h7E;
mem[16'hB6C3] = 8'hDA;
mem[16'hB6C4] = 8'hA0;
mem[16'hB6C5] = 8'hF1;
mem[16'hB6C6] = 8'h43;
mem[16'hB6C7] = 8'hAB;
mem[16'hB6C8] = 8'hFD;
mem[16'hB6C9] = 8'h65;
mem[16'hB6CA] = 8'hCB;
mem[16'hB6CB] = 8'hFF;
mem[16'hB6CC] = 8'h49;
mem[16'hB6CD] = 8'h62;
mem[16'hB6CE] = 8'hFB;
mem[16'hB6CF] = 8'h63;
mem[16'hB6D0] = 8'hD3;
mem[16'hB6D1] = 8'hB5;
mem[16'hB6D2] = 8'hAE;
mem[16'hB6D3] = 8'h8E;
mem[16'hB6D4] = 8'h18;
mem[16'hB6D5] = 8'h79;
mem[16'hB6D6] = 8'h7A;
mem[16'hB6D7] = 8'h7B;
mem[16'hB6D8] = 8'h54;
mem[16'hB6D9] = 8'h9A;
mem[16'hB6DA] = 8'hC0;
mem[16'hB6DB] = 8'hDA;
mem[16'hB6DC] = 8'h78;
mem[16'hB6DD] = 8'hD1;
mem[16'hB6DE] = 8'h82;
mem[16'hB6DF] = 8'h7D;
mem[16'hB6E0] = 8'hE5;
mem[16'hB6E1] = 8'hD5;
mem[16'hB6E2] = 8'hCB;
mem[16'hB6E3] = 8'h4F;
mem[16'hB6E4] = 8'hE1;
mem[16'hB6E5] = 8'h49;
mem[16'hB6E6] = 8'hCF;
mem[16'hB6E7] = 8'h4A;
mem[16'hB6E8] = 8'h64;
mem[16'hB6E9] = 8'h4A;
mem[16'hB6EA] = 8'hF3;
mem[16'hB6EB] = 8'h67;
mem[16'hB6EC] = 8'hAF;
mem[16'hB6ED] = 8'hF7;
mem[16'hB6EE] = 8'h22;
mem[16'hB6EF] = 8'hE3;
mem[16'hB6F0] = 8'h63;
mem[16'hB6F1] = 8'h7D;
mem[16'hB6F2] = 8'h52;
mem[16'hB6F3] = 8'hEA;
mem[16'hB6F4] = 8'hF1;
mem[16'hB6F5] = 8'hD5;
mem[16'hB6F6] = 8'h5F;
mem[16'hB6F7] = 8'h51;
mem[16'hB6F8] = 8'hD9;
mem[16'hB6F9] = 8'h35;
mem[16'hB6FA] = 8'hE1;
mem[16'hB6FB] = 8'hDA;
mem[16'hB6FC] = 8'h3D;
mem[16'hB6FD] = 8'hE6;
mem[16'hB6FE] = 8'hDF;
mem[16'hB6FF] = 8'hD3;
mem[16'hB700] = 8'h1B;
mem[16'hB701] = 8'h20;
mem[16'hB702] = 8'h3D;
mem[16'hB703] = 8'h18;
mem[16'hB704] = 8'h25;
mem[16'hB705] = 8'h01;
mem[16'hB706] = 8'h1D;
mem[16'hB707] = 8'h26;
mem[16'hB708] = 8'h1A;
mem[16'hB709] = 8'h12;
mem[16'hB70A] = 8'h04;
mem[16'hB70B] = 8'hA7;
mem[16'hB70C] = 8'h26;
mem[16'hB70D] = 8'hB7;
mem[16'hB70E] = 8'h2C;
mem[16'hB70F] = 8'hAB;
mem[16'hB710] = 8'h1C;
mem[16'hB711] = 8'h00;
mem[16'hB712] = 8'hBE;
mem[16'hB713] = 8'h16;
mem[16'hB714] = 8'h35;
mem[16'hB715] = 8'hCF;
mem[16'hB716] = 8'h0D;
mem[16'hB717] = 8'h36;
mem[16'hB718] = 8'h3D;
mem[16'hB719] = 8'h02;
mem[16'hB71A] = 8'h3B;
mem[16'hB71B] = 8'h2B;
mem[16'hB71C] = 8'h07;
mem[16'hB71D] = 8'h17;
mem[16'hB71E] = 8'hA4;
mem[16'hB71F] = 8'h0E;
mem[16'hB720] = 8'h8C;
mem[16'hB721] = 8'h27;
mem[16'hB722] = 8'h0B;
mem[16'hB723] = 8'h8E;
mem[16'hB724] = 8'hA8;
mem[16'hB725] = 8'h86;
mem[16'hB726] = 8'h3F;
mem[16'hB727] = 8'h2E;
mem[16'hB728] = 8'h83;
mem[16'hB729] = 8'h8C;
mem[16'hB72A] = 8'h87;
mem[16'hB72B] = 8'h02;
mem[16'hB72C] = 8'h87;
mem[16'hB72D] = 8'hCD;
mem[16'hB72E] = 8'hB4;
mem[16'hB72F] = 8'h34;
mem[16'hB730] = 8'h39;
mem[16'hB731] = 8'h9A;
mem[16'hB732] = 8'hB7;
mem[16'hB733] = 8'h61;
mem[16'hB734] = 8'h1D;
mem[16'hB735] = 8'h9E;
mem[16'hB736] = 8'hBA;
mem[16'hB737] = 8'h9D;
mem[16'hB738] = 8'h21;
mem[16'hB739] = 8'h28;
mem[16'hB73A] = 8'h1A;
mem[16'hB73B] = 8'h57;
mem[16'hB73C] = 8'h80;
mem[16'hB73D] = 8'h6A;
mem[16'hB73E] = 8'h5B;
mem[16'hB73F] = 8'h79;
mem[16'hB740] = 8'h3C;
mem[16'hB741] = 8'h19;
mem[16'hB742] = 8'h4E;
mem[16'hB743] = 8'hFB;
mem[16'hB744] = 8'h55;
mem[16'hB745] = 8'h65;
mem[16'hB746] = 8'h2A;
mem[16'hB747] = 8'hFB;
mem[16'hB748] = 8'h1F;
mem[16'hB749] = 8'h2C;
mem[16'hB74A] = 8'h7C;
mem[16'hB74B] = 8'h17;
mem[16'hB74C] = 8'hE9;
mem[16'hB74D] = 8'h69;
mem[16'hB74E] = 8'h32;
mem[16'hB74F] = 8'h17;
mem[16'hB750] = 8'h55;
mem[16'hB751] = 8'hEF;
mem[16'hB752] = 8'h73;
mem[16'hB753] = 8'hF7;
mem[16'hB754] = 8'h58;
mem[16'hB755] = 8'h99;
mem[16'hB756] = 8'h5A;
mem[16'hB757] = 8'hAE;
mem[16'hB758] = 8'h52;
mem[16'hB759] = 8'hE3;
mem[16'hB75A] = 8'h5F;
mem[16'hB75B] = 8'hF7;
mem[16'hB75C] = 8'h1A;
mem[16'hB75D] = 8'h74;
mem[16'hB75E] = 8'hFF;
mem[16'hB75F] = 8'h5E;
mem[16'hB760] = 8'h20;
mem[16'hB761] = 8'h0D;
mem[16'hB762] = 8'hDE;
mem[16'hB763] = 8'h34;
mem[16'hB764] = 8'h62;
mem[16'hB765] = 8'h8C;
mem[16'hB766] = 8'hC7;
mem[16'hB767] = 8'h4E;
mem[16'hB768] = 8'hC9;
mem[16'hB769] = 8'h78;
mem[16'hB76A] = 8'hC6;
mem[16'hB76B] = 8'h6B;
mem[16'hB76C] = 8'h6E;
mem[16'hB76D] = 8'h2D;
mem[16'hB76E] = 8'h02;
mem[16'hB76F] = 8'hD3;
mem[16'hB770] = 8'h27;
mem[16'hB771] = 8'hC0;
mem[16'hB772] = 8'hDE;
mem[16'hB773] = 8'h72;
mem[16'hB774] = 8'h41;
mem[16'hB775] = 8'h73;
mem[16'hB776] = 8'h25;
mem[16'hB777] = 8'h51;
mem[16'hB778] = 8'h91;
mem[16'hB779] = 8'hD8;
mem[16'hB77A] = 8'h53;
mem[16'hB77B] = 8'hDA;
mem[16'hB77C] = 8'h6D;
mem[16'hB77D] = 8'hD1;
mem[16'hB77E] = 8'h7C;
mem[16'hB77F] = 8'h7D;
mem[16'hB780] = 8'hC0;
mem[16'hB781] = 8'hED;
mem[16'hB782] = 8'h3E;
mem[16'hB783] = 8'hD4;
mem[16'hB784] = 8'h35;
mem[16'hB785] = 8'h29;
mem[16'hB786] = 8'h85;
mem[16'hB787] = 8'hB2;
mem[16'hB788] = 8'h72;
mem[16'hB789] = 8'hDA;
mem[16'hB78A] = 8'hAC;
mem[16'hB78B] = 8'h62;
mem[16'hB78C] = 8'h2D;
mem[16'hB78D] = 8'hA4;
mem[16'hB78E] = 8'h2F;
mem[16'hB78F] = 8'h9E;
mem[16'hB790] = 8'h3C;
mem[16'hB791] = 8'h8D;
mem[16'hB792] = 8'h90;
mem[16'hB793] = 8'hD3;
mem[16'hB794] = 8'hF8;
mem[16'hB795] = 8'h29;
mem[16'hB796] = 8'hC1;
mem[16'hB797] = 8'h26;
mem[16'hB798] = 8'h34;
mem[16'hB799] = 8'h84;
mem[16'hB79A] = 8'hAF;
mem[16'hB79B] = 8'h37;
mem[16'hB79C] = 8'hCF;
mem[16'hB79D] = 8'hBB;
mem[16'hB79E] = 8'h77;
mem[16'hB79F] = 8'h3E;
mem[16'hB7A0] = 8'h89;
mem[16'hB7A1] = 8'h00;
mem[16'hB7A2] = 8'h86;
mem[16'hB7A3] = 8'h1F;
mem[16'hB7A4] = 8'hB2;
mem[16'hB7A5] = 8'hAF;
mem[16'hB7A6] = 8'h1C;
mem[16'hB7A7] = 8'hA6;
mem[16'hB7A8] = 8'hE8;
mem[16'hB7A9] = 8'hC5;
mem[16'hB7AA] = 8'h16;
mem[16'hB7AB] = 8'hFC;
mem[16'hB7AC] = 8'hC9;
mem[16'hB7AD] = 8'h9A;
mem[16'hB7AE] = 8'hD2;
mem[16'hB7AF] = 8'h45;
mem[16'hB7B0] = 8'hF4;
mem[16'hB7B1] = 8'hA0;
mem[16'hB7B2] = 8'h1E;
mem[16'hB7B3] = 8'hB6;
mem[16'hB7B4] = 8'h95;
mem[16'hB7B5] = 8'h6F;
mem[16'hB7B6] = 8'hAD;
mem[16'hB7B7] = 8'h96;
mem[16'hB7B8] = 8'h9D;
mem[16'hB7B9] = 8'hA2;
mem[16'hB7BA] = 8'h9B;
mem[16'hB7BB] = 8'h8B;
mem[16'hB7BC] = 8'hA7;
mem[16'hB7BD] = 8'hBC;
mem[16'hB7BE] = 8'hFE;
mem[16'hB7BF] = 8'hD3;
mem[16'hB7C0] = 8'h7C;
mem[16'hB7C1] = 8'h96;
mem[16'hB7C2] = 8'h2B;
mem[16'hB7C3] = 8'h62;
mem[16'hB7C4] = 8'h41;
mem[16'hB7C5] = 8'h3C;
mem[16'hB7C6] = 8'hBA;
mem[16'hB7C7] = 8'h43;
mem[16'hB7C8] = 8'hE2;
mem[16'hB7C9] = 8'h73;
mem[16'hB7CA] = 8'hC0;
mem[16'hB7CB] = 8'h6D;
mem[16'hB7CC] = 8'hDD;
mem[16'hB7CD] = 8'hED;
mem[16'hB7CE] = 8'hA2;
mem[16'hB7CF] = 8'h73;
mem[16'hB7D0] = 8'h87;
mem[16'hB7D1] = 8'h77;
mem[16'hB7D2] = 8'h3B;
mem[16'hB7D3] = 8'h72;
mem[16'hB7D4] = 8'h51;
mem[16'hB7D5] = 8'hD3;
mem[16'hB7D6] = 8'hAA;
mem[16'hB7D7] = 8'h63;
mem[16'hB7D8] = 8'hD2;
mem[16'hB7D9] = 8'h63;
mem[16'hB7DA] = 8'hCB;
mem[16'hB7DB] = 8'h77;
mem[16'hB7DC] = 8'hD9;
mem[16'hB7DD] = 8'h81;
mem[16'hB7DE] = 8'h6E;
mem[16'hB7DF] = 8'hCE;
mem[16'hB7E0] = 8'h4C;
mem[16'hB7E1] = 8'hE7;
mem[16'hB7E2] = 8'h8B;
mem[16'hB7E3] = 8'h4F;
mem[16'hB7E4] = 8'h98;
mem[16'hB7E5] = 8'h4A;
mem[16'hB7E6] = 8'h06;
mem[16'hB7E7] = 8'h7B;
mem[16'hB7E8] = 8'hF3;
mem[16'hB7E9] = 8'h8C;
mem[16'hB7EA] = 8'hB9;
mem[16'hB7EB] = 8'hB7;
mem[16'hB7EC] = 8'h4E;
mem[16'hB7ED] = 8'h0D;
mem[16'hB7EE] = 8'h5F;
mem[16'hB7EF] = 8'hF4;
mem[16'hB7F0] = 8'hF5;
mem[16'hB7F1] = 8'h49;
mem[16'hB7F2] = 8'hD3;
mem[16'hB7F3] = 8'h57;
mem[16'hB7F4] = 8'hF8;
mem[16'hB7F5] = 8'h39;
mem[16'hB7F6] = 8'hF3;
mem[16'hB7F7] = 8'h48;
mem[16'hB7F8] = 8'hD9;
mem[16'hB7F9] = 8'h5D;
mem[16'hB7FA] = 8'hF6;
mem[16'hB7FB] = 8'h37;
mem[16'hB7FC] = 8'h50;
mem[16'hB7FD] = 8'h51;
mem[16'hB7FE] = 8'h52;
mem[16'hB7FF] = 8'h53;
mem[16'hB800] = 8'h09;
mem[16'hB801] = 8'h97;
mem[16'hB802] = 8'hEB;
mem[16'hB803] = 8'h95;
mem[16'hB804] = 8'h25;
mem[16'hB805] = 8'hA0;
mem[16'hB806] = 8'h0A;
mem[16'hB807] = 8'h2E;
mem[16'hB808] = 8'hB0;
mem[16'hB809] = 8'h0C;
mem[16'hB80A] = 8'hAA;
mem[16'hB80B] = 8'h22;
mem[16'hB80C] = 8'hB5;
mem[16'hB80D] = 8'h08;
mem[16'hB80E] = 8'h5A;
mem[16'hB80F] = 8'h26;
mem[16'hB810] = 8'hAA;
mem[16'hB811] = 8'h9D;
mem[16'hB812] = 8'hC4;
mem[16'hB813] = 8'h0B;
mem[16'hB814] = 8'h18;
mem[16'hB815] = 8'hB9;
mem[16'hB816] = 8'h3E;
mem[16'hB817] = 8'hB3;
mem[16'hB818] = 8'h1D;
mem[16'hB819] = 8'hB1;
mem[16'hB81A] = 8'h33;
mem[16'hB81B] = 8'hBE;
mem[16'hB81C] = 8'h19;
mem[16'hB81D] = 8'h11;
mem[16'hB81E] = 8'h23;
mem[16'hB81F] = 8'hBB;
mem[16'hB820] = 8'h44;
mem[16'hB821] = 8'h5D;
mem[16'hB822] = 8'h75;
mem[16'hB823] = 8'h69;
mem[16'hB824] = 8'h81;
mem[16'hB825] = 8'h2C;
mem[16'hB826] = 8'h83;
mem[16'hB827] = 8'h42;
mem[16'hB828] = 8'h8C;
mem[16'hB829] = 8'h15;
mem[16'hB82A] = 8'h77;
mem[16'hB82B] = 8'h27;
mem[16'hB82C] = 8'hA7;
mem[16'hB82D] = 8'h38;
mem[16'hB82E] = 8'h56;
mem[16'hB82F] = 8'h37;
mem[16'hB830] = 8'h05;
mem[16'hB831] = 8'h9D;
mem[16'hB832] = 8'h9A;
mem[16'hB833] = 8'h17;
mem[16'hB834] = 8'h88;
mem[16'hB835] = 8'h6E;
mem[16'hB836] = 8'hBA;
mem[16'hB837] = 8'h9F;
mem[16'hB838] = 8'h2F;
mem[16'hB839] = 8'h38;
mem[16'hB83A] = 8'h86;
mem[16'hB83B] = 8'h37;
mem[16'hB83C] = 8'hB9;
mem[16'hB83D] = 8'h3B;
mem[16'hB83E] = 8'hD8;
mem[16'hB83F] = 8'h9A;
mem[16'hB840] = 8'h64;
mem[16'hB841] = 8'hC0;
mem[16'hB842] = 8'hFE;
mem[16'hB843] = 8'h4F;
mem[16'hB844] = 8'h38;
mem[16'hB845] = 8'hB5;
mem[16'hB846] = 8'h43;
mem[16'hB847] = 8'hEA;
mem[16'hB848] = 8'h61;
mem[16'hB849] = 8'hEC;
mem[16'hB84A] = 8'h4B;
mem[16'hB84B] = 8'h64;
mem[16'hB84C] = 8'h20;
mem[16'hB84D] = 8'h6C;
mem[16'hB84E] = 8'hFE;
mem[16'hB84F] = 8'h43;
mem[16'hB850] = 8'h51;
mem[16'hB851] = 8'h7E;
mem[16'hB852] = 8'h3E;
mem[16'hB853] = 8'h72;
mem[16'hB854] = 8'hE3;
mem[16'hB855] = 8'h59;
mem[16'hB856] = 8'h53;
mem[16'hB857] = 8'h04;
mem[16'hB858] = 8'h65;
mem[16'hB859] = 8'hFD;
mem[16'hB85A] = 8'h27;
mem[16'hB85B] = 8'hFF;
mem[16'hB85C] = 8'h20;
mem[16'hB85D] = 8'hFD;
mem[16'hB85E] = 8'h5B;
mem[16'hB85F] = 8'hF3;
mem[16'hB860] = 8'h5D;
mem[16'hB861] = 8'hC5;
mem[16'hB862] = 8'h06;
mem[16'hB863] = 8'h07;
mem[16'hB864] = 8'h18;
mem[16'hB865] = 8'h33;
mem[16'hB866] = 8'h1B;
mem[16'hB867] = 8'hC3;
mem[16'hB868] = 8'h34;
mem[16'hB869] = 8'hC8;
mem[16'hB86A] = 8'h63;
mem[16'hB86B] = 8'hCE;
mem[16'hB86C] = 8'h09;
mem[16'hB86D] = 8'h01;
mem[16'hB86E] = 8'h52;
mem[16'hB86F] = 8'hF1;
mem[16'hB870] = 8'h75;
mem[16'hB871] = 8'h1D;
mem[16'hB872] = 8'h53;
mem[16'hB873] = 8'hC6;
mem[16'hB874] = 8'h78;
mem[16'hB875] = 8'hE9;
mem[16'hB876] = 8'hD1;
mem[16'hB877] = 8'h7E;
mem[16'hB878] = 8'hDD;
mem[16'hB879] = 8'h1C;
mem[16'hB87A] = 8'h06;
mem[16'hB87B] = 8'h47;
mem[16'hB87C] = 8'hD5;
mem[16'hB87D] = 8'h78;
mem[16'hB87E] = 8'hD2;
mem[16'hB87F] = 8'h5E;
mem[16'hB880] = 8'h35;
mem[16'hB881] = 8'h8D;
mem[16'hB882] = 8'hC8;
mem[16'hB883] = 8'h26;
mem[16'hB884] = 8'hD8;
mem[16'hB885] = 8'h08;
mem[16'hB886] = 8'h8F;
mem[16'hB887] = 8'h22;
mem[16'hB888] = 8'hED;
mem[16'hB889] = 8'h85;
mem[16'hB88A] = 8'hD6;
mem[16'hB88B] = 8'hD1;
mem[16'hB88C] = 8'hE9;
mem[16'hB88D] = 8'h25;
mem[16'hB88E] = 8'hB2;
mem[16'hB88F] = 8'hE5;
mem[16'hB890] = 8'hF5;
mem[16'hB891] = 8'h35;
mem[16'hB892] = 8'hAE;
mem[16'hB893] = 8'hD1;
mem[16'hB894] = 8'hF1;
mem[16'hB895] = 8'h91;
mem[16'hB896] = 8'hAA;
mem[16'hB897] = 8'h85;
mem[16'hB898] = 8'hFD;
mem[16'hB899] = 8'hF5;
mem[16'hB89A] = 8'hA6;
mem[16'hB89B] = 8'hD1;
mem[16'hB89C] = 8'hF9;
mem[16'hB89D] = 8'hF1;
mem[16'hB89E] = 8'hC2;
mem[16'hB89F] = 8'hD1;
mem[16'hB8A0] = 8'hDC;
mem[16'hB8A1] = 8'hB9;
mem[16'hB8A2] = 8'hA7;
mem[16'hB8A3] = 8'h06;
mem[16'hB8A4] = 8'h44;
mem[16'hB8A5] = 8'h09;
mem[16'hB8A6] = 8'hB1;
mem[16'hB8A7] = 8'h47;
mem[16'hB8A8] = 8'hE4;
mem[16'hB8A9] = 8'hB7;
mem[16'hB8AA] = 8'h06;
mem[16'hB8AB] = 8'h07;
mem[16'hB8AC] = 8'h00;
mem[16'hB8AD] = 8'h01;
mem[16'hB8AE] = 8'h02;
mem[16'hB8AF] = 8'h03;
mem[16'hB8B0] = 8'hB5;
mem[16'hB8B1] = 8'h91;
mem[16'hB8B2] = 8'h1B;
mem[16'hB8B3] = 8'h15;
mem[16'hB8B4] = 8'h95;
mem[16'hB8B5] = 8'h83;
mem[16'hB8B6] = 8'hA3;
mem[16'hB8B7] = 8'h96;
mem[16'hB8B8] = 8'hA5;
mem[16'hB8B9] = 8'hAC;
mem[16'hB8BA] = 8'h9B;
mem[16'hB8BB] = 8'hDE;
mem[16'hB8BC] = 8'hA9;
mem[16'hB8BD] = 8'h9C;
mem[16'hB8BE] = 8'hF2;
mem[16'hB8BF] = 8'hAA;
mem[16'hB8C0] = 8'hE1;
mem[16'hB8C1] = 8'h9A;
mem[16'hB8C2] = 8'hD7;
mem[16'hB8C3] = 8'hE2;
mem[16'hB8C4] = 8'h67;
mem[16'hB8C5] = 8'hD3;
mem[16'hB8C6] = 8'hC3;
mem[16'hB8C7] = 8'hE6;
mem[16'hB8C8] = 8'h61;
mem[16'hB8C9] = 8'h6F;
mem[16'hB8CA] = 8'hEB;
mem[16'hB8CB] = 8'hF0;
mem[16'hB8CC] = 8'hD9;
mem[16'hB8CD] = 8'hEC;
mem[16'hB8CE] = 8'hCC;
mem[16'hB8CF] = 8'hDA;
mem[16'hB8D0] = 8'hF1;
mem[16'hB8D1] = 8'hBB;
mem[16'hB8D2] = 8'hC7;
mem[16'hB8D3] = 8'hF2;
mem[16'hB8D4] = 8'hA5;
mem[16'hB8D5] = 8'hC0;
mem[16'hB8D6] = 8'hF7;
mem[16'hB8D7] = 8'h8F;
mem[16'hB8D8] = 8'hCD;
mem[16'hB8D9] = 8'hF8;
mem[16'hB8DA] = 8'h7A;
mem[16'hB8DB] = 8'hCD;
mem[16'hB8DC] = 8'hD2;
mem[16'hB8DD] = 8'h71;
mem[16'hB8DE] = 8'hF4;
mem[16'hB8DF] = 8'h65;
mem[16'hB8E0] = 8'hF1;
mem[16'hB8E1] = 8'h4D;
mem[16'hB8E2] = 8'hE7;
mem[16'hB8E3] = 8'hC2;
mem[16'hB8E4] = 8'hC7;
mem[16'hB8E5] = 8'hF0;
mem[16'hB8E6] = 8'hC7;
mem[16'hB8E7] = 8'hE9;
mem[16'hB8E8] = 8'hFD;
mem[16'hB8E9] = 8'hC8;
mem[16'hB8EA] = 8'hFF;
mem[16'hB8EB] = 8'hFE;
mem[16'hB8EC] = 8'hCD;
mem[16'hB8ED] = 8'h90;
mem[16'hB8EE] = 8'hFB;
mem[16'hB8EF] = 8'hCE;
mem[16'hB8F0] = 8'h84;
mem[16'hB8F1] = 8'hE4;
mem[16'hB8F2] = 8'hE3;
mem[16'hB8F3] = 8'h5F;
mem[16'hB8F4] = 8'hF2;
mem[16'hB8F5] = 8'hDC;
mem[16'hB8F6] = 8'h5B;
mem[16'hB8F7] = 8'h7B;
mem[16'hB8F8] = 8'h5B;
mem[16'hB8F9] = 8'hE0;
mem[16'hB8FA] = 8'hF6;
mem[16'hB8FB] = 8'h68;
mem[16'hB8FC] = 8'h1C;
mem[16'hB8FD] = 8'h58;
mem[16'hB8FE] = 8'hE7;
mem[16'hB8FF] = 8'h53;
mem[16'hB900] = 8'hE0;
mem[16'hB901] = 8'h35;
mem[16'hB902] = 8'h14;
mem[16'hB903] = 8'h8F;
mem[16'hB904] = 8'h18;
mem[16'hB905] = 8'h11;
mem[16'hB906] = 8'h8A;
mem[16'hB907] = 8'h1F;
mem[16'hB908] = 8'h1E;
mem[16'hB909] = 8'h03;
mem[16'hB90A] = 8'hAC;
mem[16'hB90B] = 8'h07;
mem[16'hB90C] = 8'hA4;
mem[16'hB90D] = 8'h08;
mem[16'hB90E] = 8'h5D;
mem[16'hB90F] = 8'h3E;
mem[16'hB910] = 8'h33;
mem[16'hB911] = 8'h7D;
mem[16'hB912] = 8'h63;
mem[16'hB913] = 8'h33;
mem[16'hB914] = 8'h78;
mem[16'hB915] = 8'h53;
mem[16'hB916] = 8'h7F;
mem[16'hB917] = 8'hAD;
mem[16'hB918] = 8'h94;
mem[16'hB919] = 8'hE2;
mem[16'hB91A] = 8'h0C;
mem[16'hB91B] = 8'h72;
mem[16'hB91C] = 8'hA0;
mem[16'hB91D] = 8'h2C;
mem[16'hB91E] = 8'h3F;
mem[16'hB91F] = 8'h73;
mem[16'hB920] = 8'h51;
mem[16'hB921] = 8'h01;
mem[16'hB922] = 8'h4E;
mem[16'hB923] = 8'h07;
mem[16'hB924] = 8'h58;
mem[16'hB925] = 8'h7B;
mem[16'hB926] = 8'hAA;
mem[16'hB927] = 8'hD3;
mem[16'hB928] = 8'h3E;
mem[16'hB929] = 8'h2C;
mem[16'hB92A] = 8'h11;
mem[16'hB92B] = 8'h1A;
mem[16'hB92C] = 8'h0D;
mem[16'hB92D] = 8'h41;
mem[16'hB92E] = 8'h5F;
mem[16'hB92F] = 8'h0F;
mem[16'hB930] = 8'h5C;
mem[16'hB931] = 8'h33;
mem[16'hB932] = 8'h88;
mem[16'hB933] = 8'h9F;
mem[16'hB934] = 8'h25;
mem[16'hB935] = 8'h99;
mem[16'hB936] = 8'h31;
mem[16'hB937] = 8'h3D;
mem[16'hB938] = 8'h9E;
mem[16'hB939] = 8'hB5;
mem[16'hB93A] = 8'hCD;
mem[16'hB93B] = 8'h2D;
mem[16'hB93C] = 8'h0D;
mem[16'hB93D] = 8'h1C;
mem[16'hB93E] = 8'h52;
mem[16'hB93F] = 8'h4E;
mem[16'hB940] = 8'h60;
mem[16'hB941] = 8'h2D;
mem[16'hB942] = 8'h47;
mem[16'hB943] = 8'h05;
mem[16'hB944] = 8'hC8;
mem[16'hB945] = 8'hB1;
mem[16'hB946] = 8'h50;
mem[16'hB947] = 8'h76;
mem[16'hB948] = 8'h69;
mem[16'hB949] = 8'h25;
mem[16'hB94A] = 8'h3B;
mem[16'hB94B] = 8'h6B;
mem[16'hB94C] = 8'h20;
mem[16'hB94D] = 8'hC1;
mem[16'hB94E] = 8'hB1;
mem[16'hB94F] = 8'h5A;
mem[16'hB950] = 8'h2C;
mem[16'hB951] = 8'h4A;
mem[16'hB952] = 8'h9E;
mem[16'hB953] = 8'h5F;
mem[16'hB954] = 8'hF3;
mem[16'hB955] = 8'h50;
mem[16'hB956] = 8'h05;
mem[16'hB957] = 8'hB7;
mem[16'hB958] = 8'hAA;
mem[16'hB959] = 8'h4C;
mem[16'hB95A] = 8'hD6;
mem[16'hB95B] = 8'hAD;
mem[16'hB95C] = 8'h4A;
mem[16'hB95D] = 8'h1B;
mem[16'hB95E] = 8'hBA;
mem[16'hB95F] = 8'h9B;
mem[16'hB960] = 8'h09;
mem[16'hB961] = 8'hCD;
mem[16'hB962] = 8'h53;
mem[16'hB963] = 8'h42;
mem[16'hB964] = 8'h08;
mem[16'hB965] = 8'h14;
mem[16'hB966] = 8'h46;
mem[16'hB967] = 8'h0B;
mem[16'hB968] = 8'h4C;
mem[16'hB969] = 8'h15;
mem[16'hB96A] = 8'h29;
mem[16'hB96B] = 8'h2D;
mem[16'hB96C] = 8'h6D;
mem[16'hB96D] = 8'h4E;
mem[16'hB96E] = 8'h7B;
mem[16'hB96F] = 8'h63;
mem[16'hB970] = 8'h89;
mem[16'hB971] = 8'h7B;
mem[16'hB972] = 8'hD4;
mem[16'hB973] = 8'h52;
mem[16'hB974] = 8'hA0;
mem[16'hB975] = 8'h60;
mem[16'hB976] = 8'h63;
mem[16'hB977] = 8'hDB;
mem[16'hB978] = 8'hF4;
mem[16'hB979] = 8'h58;
mem[16'hB97A] = 8'h6B;
mem[16'hB97B] = 8'h6E;
mem[16'hB97C] = 8'h79;
mem[16'hB97D] = 8'h4B;
mem[16'hB97E] = 8'h38;
mem[16'hB97F] = 8'h4E;
mem[16'hB980] = 8'hA1;
mem[16'hB981] = 8'hED;
mem[16'hB982] = 8'hF3;
mem[16'hB983] = 8'hA3;
mem[16'hB984] = 8'hE8;
mem[16'hB985] = 8'h87;
mem[16'hB986] = 8'h3C;
mem[16'hB987] = 8'h2B;
mem[16'hB988] = 8'h8D;
mem[16'hB989] = 8'h25;
mem[16'hB98A] = 8'hCC;
mem[16'hB98B] = 8'hA2;
mem[16'hB98C] = 8'h2D;
mem[16'hB98D] = 8'h9F;
mem[16'hB98E] = 8'h88;
mem[16'hB98F] = 8'h03;
mem[16'hB990] = 8'hD6;
mem[16'hB991] = 8'hF8;
mem[16'hB992] = 8'h2E;
mem[16'hB993] = 8'h82;
mem[16'hB994] = 8'h38;
mem[16'hB995] = 8'h95;
mem[16'hB996] = 8'hB7;
mem[16'hB997] = 8'hB6;
mem[16'hB998] = 8'hF4;
mem[16'hB999] = 8'hF8;
mem[16'hB99A] = 8'hBA;
mem[16'hB99B] = 8'hF7;
mem[16'hB99C] = 8'h75;
mem[16'hB99D] = 8'h3C;
mem[16'hB99E] = 8'hB7;
mem[16'hB99F] = 8'h3E;
mem[16'hB9A0] = 8'hB5;
mem[16'hB9A1] = 8'h5B;
mem[16'hB9A2] = 8'h2E;
mem[16'hB9A3] = 8'h26;
mem[16'hB9A4] = 8'h07;
mem[16'hB9A5] = 8'h14;
mem[16'hB9A6] = 8'h0A;
mem[16'hB9A7] = 8'hA6;
mem[16'hB9A8] = 8'hAE;
mem[16'hB9A9] = 8'hB8;
mem[16'hB9AA] = 8'h06;
mem[16'hB9AB] = 8'hA9;
mem[16'hB9AC] = 8'hEA;
mem[16'hB9AD] = 8'h8C;
mem[16'hB9AE] = 8'h8F;
mem[16'hB9AF] = 8'hC3;
mem[16'hB9B0] = 8'hD1;
mem[16'hB9B1] = 8'h91;
mem[16'hB9B2] = 8'hDE;
mem[16'hB9B3] = 8'h5A;
mem[16'hB9B4] = 8'h15;
mem[16'hB9B5] = 8'h9C;
mem[16'hB9B6] = 8'h17;
mem[16'hB9B7] = 8'hA2;
mem[16'hB9B8] = 8'h42;
mem[16'hB9B9] = 8'h35;
mem[16'hB9BA] = 8'h3F;
mem[16'hB9BB] = 8'hE7;
mem[16'hB9BC] = 8'hB2;
mem[16'hB9BD] = 8'h11;
mem[16'hB9BE] = 8'h0F;
mem[16'hB9BF] = 8'h13;
mem[16'hB9C0] = 8'hC3;
mem[16'hB9C1] = 8'hC7;
mem[16'hB9C2] = 8'hD3;
mem[16'hB9C3] = 8'h6F;
mem[16'hB9C4] = 8'hD8;
mem[16'hB9C5] = 8'hE4;
mem[16'hB9C6] = 8'hE7;
mem[16'hB9C7] = 8'hAB;
mem[16'hB9C8] = 8'hA9;
mem[16'hB9C9] = 8'hE9;
mem[16'hB9CA] = 8'hA6;
mem[16'hB9CB] = 8'h22;
mem[16'hB9CC] = 8'h6D;
mem[16'hB9CD] = 8'hE4;
mem[16'hB9CE] = 8'h6F;
mem[16'hB9CF] = 8'hDD;
mem[16'hB9D0] = 8'h7C;
mem[16'hB9D1] = 8'h5D;
mem[16'hB9D2] = 8'hC3;
mem[16'hB9D3] = 8'h7F;
mem[16'hB9D4] = 8'hC9;
mem[16'hB9D5] = 8'hF1;
mem[16'hB9D6] = 8'hC4;
mem[16'hB9D7] = 8'h7B;
mem[16'hB9D8] = 8'h54;
mem[16'hB9D9] = 8'hFB;
mem[16'hB9DA] = 8'hCB;
mem[16'hB9DB] = 8'hCE;
mem[16'hB9DC] = 8'hFD;
mem[16'hB9DD] = 8'hFC;
mem[16'hB9DE] = 8'hB2;
mem[16'hB9DF] = 8'hBE;
mem[16'hB9E0] = 8'hC0;
mem[16'hB9E1] = 8'h8D;
mem[16'hB9E2] = 8'h0B;
mem[16'hB9E3] = 8'h42;
mem[16'hB9E4] = 8'hCD;
mem[16'hB9E5] = 8'h44;
mem[16'hB9E6] = 8'h8A;
mem[16'hB9E7] = 8'h4B;
mem[16'hB9E8] = 8'h54;
mem[16'hB9E9] = 8'hE6;
mem[16'hB9EA] = 8'hA0;
mem[16'hB9EB] = 8'h51;
mem[16'hB9EC] = 8'hE6;
mem[16'hB9ED] = 8'h57;
mem[16'hB9EE] = 8'hFF;
mem[16'hB9EF] = 8'h43;
mem[16'hB9F0] = 8'hF5;
mem[16'hB9F1] = 8'hFD;
mem[16'hB9F2] = 8'hC5;
mem[16'hB9F3] = 8'hD3;
mem[16'hB9F4] = 8'hD5;
mem[16'hB9F5] = 8'h99;
mem[16'hB9F6] = 8'h96;
mem[16'hB9F7] = 8'hD7;
mem[16'hB9F8] = 8'h94;
mem[16'hB9F9] = 8'hD8;
mem[16'hB9FA] = 8'hD9;
mem[16'hB9FB] = 8'hEE;
mem[16'hB9FC] = 8'hDD;
mem[16'hB9FD] = 8'hF3;
mem[16'hB9FE] = 8'hEB;
mem[16'hB9FF] = 8'hDE;
mem[16'hBA00] = 8'h15;
mem[16'hBA01] = 8'h14;
mem[16'hBA02] = 8'h23;
mem[16'hBA03] = 8'h7E;
mem[16'hBA04] = 8'h11;
mem[16'hBA05] = 8'h01;
mem[16'hBA06] = 8'h07;
mem[16'hBA07] = 8'hA6;
mem[16'hBA08] = 8'hA4;
mem[16'hBA09] = 8'hAC;
mem[16'hBA0A] = 8'h0C;
mem[16'hBA0B] = 8'h2A;
mem[16'hBA0C] = 8'h2D;
mem[16'hBA0D] = 8'h61;
mem[16'hBA0E] = 8'h6F;
mem[16'hBA0F] = 8'h2F;
mem[16'hBA10] = 8'h7C;
mem[16'hBA11] = 8'h31;
mem[16'hBA12] = 8'h66;
mem[16'hBA13] = 8'h06;
mem[16'hBA14] = 8'h1D;
mem[16'hBA15] = 8'hB4;
mem[16'hBA16] = 8'hF0;
mem[16'hBA17] = 8'hB2;
mem[16'hBA18] = 8'h1E;
mem[16'hBA19] = 8'h13;
mem[16'hBA1A] = 8'hBC;
mem[16'hBA1B] = 8'hFF;
mem[16'hBA1C] = 8'hD8;
mem[16'hBA1D] = 8'h5B;
mem[16'hBA1E] = 8'h2F;
mem[16'hBA1F] = 8'h3E;
mem[16'hBA20] = 8'h4C;
mem[16'hBA21] = 8'h50;
mem[16'hBA22] = 8'h02;
mem[16'hBA23] = 8'h4F;
mem[16'hBA24] = 8'hA8;
mem[16'hBA25] = 8'hDE;
mem[16'hBA26] = 8'h30;
mem[16'hBA27] = 8'h16;
mem[16'hBA28] = 8'h09;
mem[16'hBA29] = 8'h45;
mem[16'hBA2A] = 8'h5B;
mem[16'hBA2B] = 8'h0B;
mem[16'hBA2C] = 8'h40;
mem[16'hBA2D] = 8'hA1;
mem[16'hBA2E] = 8'hD5;
mem[16'hBA2F] = 8'h39;
mem[16'hBA30] = 8'h01;
mem[16'hBA31] = 8'h10;
mem[16'hBA32] = 8'h5E;
mem[16'hBA33] = 8'h42;
mem[16'hBA34] = 8'h16;
mem[16'hBA35] = 8'h59;
mem[16'hBA36] = 8'h3C;
mem[16'hBA37] = 8'h8D;
mem[16'hBA38] = 8'h64;
mem[16'hBA39] = 8'h87;
mem[16'hBA3A] = 8'h2B;
mem[16'hBA3B] = 8'h97;
mem[16'hBA3C] = 8'h3A;
mem[16'hBA3D] = 8'h54;
mem[16'hBA3E] = 8'h92;
mem[16'hBA3F] = 8'h63;
mem[16'hBA40] = 8'hE5;
mem[16'hBA41] = 8'h68;
mem[16'hBA42] = 8'hEF;
mem[16'hBA43] = 8'h26;
mem[16'hBA44] = 8'h17;
mem[16'hBA45] = 8'h19;
mem[16'hBA46] = 8'hEF;
mem[16'hBA47] = 8'hCB;
mem[16'hBA48] = 8'hEB;
mem[16'hBA49] = 8'h50;
mem[16'hBA4A] = 8'h4F;
mem[16'hBA4B] = 8'hE6;
mem[16'hBA4C] = 8'hE8;
mem[16'hBA4D] = 8'h47;
mem[16'hBA4E] = 8'hE8;
mem[16'hBA4F] = 8'h5E;
mem[16'hBA50] = 8'h71;
mem[16'hBA51] = 8'h3D;
mem[16'hBA52] = 8'h43;
mem[16'hBA53] = 8'h71;
mem[16'hBA54] = 8'h38;
mem[16'hBA55] = 8'hD1;
mem[16'hBA56] = 8'h9A;
mem[16'hBA57] = 8'h11;
mem[16'hBA58] = 8'hBC;
mem[16'hBA59] = 8'h9D;
mem[16'hBA5A] = 8'h1C;
mem[16'hBA5B] = 8'h97;
mem[16'hBA5C] = 8'hD0;
mem[16'hBA5D] = 8'h41;
mem[16'hBA5E] = 8'h4A;
mem[16'hBA5F] = 8'h5A;
mem[16'hBA60] = 8'h42;
mem[16'hBA61] = 8'h40;
mem[16'hBA62] = 8'hFA;
mem[16'hBA63] = 8'h75;
mem[16'hBA64] = 8'h6D;
mem[16'hBA65] = 8'hCE;
mem[16'hBA66] = 8'hC3;
mem[16'hBA67] = 8'hCA;
mem[16'hBA68] = 8'h41;
mem[16'hBA69] = 8'hC2;
mem[16'hBA6A] = 8'h16;
mem[16'hBA6B] = 8'hC1;
mem[16'hBA6C] = 8'h65;
mem[16'hBA6D] = 8'hC6;
mem[16'hBA6E] = 8'hEB;
mem[16'hBA6F] = 8'h3D;
mem[16'hBA70] = 8'h59;
mem[16'hBA71] = 8'hDA;
mem[16'hBA72] = 8'h77;
mem[16'hBA73] = 8'hDC;
mem[16'hBA74] = 8'h5D;
mem[16'hBA75] = 8'hC3;
mem[16'hBA76] = 8'hFA;
mem[16'hBA77] = 8'hDD;
mem[16'hBA78] = 8'h61;
mem[16'hBA79] = 8'h68;
mem[16'hBA7A] = 8'h5A;
mem[16'hBA7B] = 8'h17;
mem[16'hBA7C] = 8'hC0;
mem[16'hBA7D] = 8'h2A;
mem[16'hBA7E] = 8'h1B;
mem[16'hBA7F] = 8'h39;
mem[16'hBA80] = 8'hFC;
mem[16'hBA81] = 8'hDD;
mem[16'hBA82] = 8'h87;
mem[16'hBA83] = 8'hD0;
mem[16'hBA84] = 8'hF5;
mem[16'hBA85] = 8'hA4;
mem[16'hBA86] = 8'hEA;
mem[16'hBA87] = 8'hB6;
mem[16'hBA88] = 8'hAB;
mem[16'hBA89] = 8'hE5;
mem[16'hBA8A] = 8'hFB;
mem[16'hBA8B] = 8'hAB;
mem[16'hBA8C] = 8'hE0;
mem[16'hBA8D] = 8'h85;
mem[16'hBA8E] = 8'h38;
mem[16'hBA8F] = 8'h03;
mem[16'hBA90] = 8'h67;
mem[16'hBA91] = 8'h87;
mem[16'hBA92] = 8'h1E;
mem[16'hBA93] = 8'h61;
mem[16'hBA94] = 8'h81;
mem[16'hBA95] = 8'hE9;
mem[16'hBA96] = 8'hEF;
mem[16'hBA97] = 8'h5B;
mem[16'hBA98] = 8'h14;
mem[16'hBA99] = 8'h69;
mem[16'hBA9A] = 8'h8C;
mem[16'hBA9B] = 8'h9A;
mem[16'hBA9C] = 8'h38;
mem[16'hBA9D] = 8'h91;
mem[16'hBA9E] = 8'hFB;
mem[16'hBA9F] = 8'h22;
mem[16'hBAA0] = 8'hDC;
mem[16'hBAA1] = 8'h1C;
mem[16'hBAA2] = 8'hA7;
mem[16'hBAA3] = 8'h0F;
mem[16'hBAA4] = 8'h8D;
mem[16'hBAA5] = 8'h08;
mem[16'hBAA6] = 8'h87;
mem[16'hBAA7] = 8'h03;
mem[16'hBAA8] = 8'hA4;
mem[16'hBAA9] = 8'hAC;
mem[16'hBAAA] = 8'h9E;
mem[16'hBAAB] = 8'h82;
mem[16'hBAAC] = 8'h00;
mem[16'hBAAD] = 8'h21;
mem[16'hBAAE] = 8'h0D;
mem[16'hBAAF] = 8'hB6;
mem[16'hBAB0] = 8'h3C;
mem[16'hBAB1] = 8'h41;
mem[16'hBAB2] = 8'hA4;
mem[16'hBAB3] = 8'h7F;
mem[16'hBAB4] = 8'hBE;
mem[16'hBAB5] = 8'h13;
mem[16'hBAB6] = 8'hA7;
mem[16'hBAB7] = 8'h96;
mem[16'hBAB8] = 8'hD4;
mem[16'hBAB9] = 8'hA8;
mem[16'hBABA] = 8'h98;
mem[16'hBABB] = 8'hD7;
mem[16'hBABC] = 8'h00;
mem[16'hBABD] = 8'h19;
mem[16'hBABE] = 8'hBB;
mem[16'hBABF] = 8'h03;
mem[16'hBAC0] = 8'hE1;
mem[16'hBAC1] = 8'h65;
mem[16'hBAC2] = 8'hCE;
mem[16'hBAC3] = 8'h07;
mem[16'hBAC4] = 8'h00;
mem[16'hBAC5] = 8'h09;
mem[16'hBAC6] = 8'hCE;
mem[16'hBAC7] = 8'h70;
mem[16'hBAC8] = 8'hF9;
mem[16'hBAC9] = 8'hEA;
mem[16'hBACA] = 8'hA6;
mem[16'hBACB] = 8'hBA;
mem[16'hBACC] = 8'hEC;
mem[16'hBACD] = 8'hA1;
mem[16'hBACE] = 8'hA4;
mem[16'hBACF] = 8'h6B;
mem[16'hBAD0] = 8'hAC;
mem[16'hBAD1] = 8'h81;
mem[16'hBAD2] = 8'hF6;
mem[16'hBAD3] = 8'hAF;
mem[16'hBAD4] = 8'h81;
mem[16'hBAD5] = 8'hC4;
mem[16'hBAD6] = 8'hF7;
mem[16'hBAD7] = 8'hBB;
mem[16'hBAD8] = 8'hC9;
mem[16'hBAD9] = 8'hFB;
mem[16'hBADA] = 8'hB6;
mem[16'hBADB] = 8'hDE;
mem[16'hBADC] = 8'hFC;
mem[16'hBADD] = 8'hFC;
mem[16'hBADE] = 8'h46;
mem[16'hBADF] = 8'hC9;
mem[16'hBAE0] = 8'h2C;
mem[16'hBAE1] = 8'h4D;
mem[16'hBAE2] = 8'h4E;
mem[16'hBAE3] = 8'h4F;
mem[16'hBAE4] = 8'h48;
mem[16'hBAE5] = 8'h49;
mem[16'hBAE6] = 8'h4A;
mem[16'hBAE7] = 8'h4B;
mem[16'hBAE8] = 8'h44;
mem[16'hBAE9] = 8'h45;
mem[16'hBAEA] = 8'h46;
mem[16'hBAEB] = 8'h47;
mem[16'hBAEC] = 8'h40;
mem[16'hBAED] = 8'h41;
mem[16'hBAEE] = 8'h42;
mem[16'hBAEF] = 8'h43;
mem[16'hBAF0] = 8'h5C;
mem[16'hBAF1] = 8'h5D;
mem[16'hBAF2] = 8'h5E;
mem[16'hBAF3] = 8'h5F;
mem[16'hBAF4] = 8'h58;
mem[16'hBAF5] = 8'h59;
mem[16'hBAF6] = 8'h5A;
mem[16'hBAF7] = 8'h5B;
mem[16'hBAF8] = 8'h54;
mem[16'hBAF9] = 8'h55;
mem[16'hBAFA] = 8'h56;
mem[16'hBAFB] = 8'h57;
mem[16'hBAFC] = 8'h50;
mem[16'hBAFD] = 8'h51;
mem[16'hBAFE] = 8'h52;
mem[16'hBAFF] = 8'h53;
mem[16'hBB00] = 8'hE0;
mem[16'hBB01] = 8'hA5;
mem[16'hBB02] = 8'h15;
mem[16'hBB03] = 8'h8F;
mem[16'hBB04] = 8'hE4;
mem[16'hBB05] = 8'hE4;
mem[16'hBB06] = 8'h14;
mem[16'hBB07] = 8'h02;
mem[16'hBB08] = 8'h6D;
mem[16'hBB09] = 8'hAF;
mem[16'hBB0A] = 8'h36;
mem[16'hBB0B] = 8'hA0;
mem[16'hBB0C] = 8'h09;
mem[16'hBB0D] = 8'hA8;
mem[16'hBB0E] = 8'h2F;
mem[16'hBB0F] = 8'hAB;
mem[16'hBB10] = 8'h1C;
mem[16'hBB11] = 8'hDD;
mem[16'hBB12] = 8'hCB;
mem[16'hBB13] = 8'h1D;
mem[16'hBB14] = 8'hB8;
mem[16'hBB15] = 8'h3F;
mem[16'hBB16] = 8'hBC;
mem[16'hBB17] = 8'h35;
mem[16'hBB18] = 8'hBC;
mem[16'hBB19] = 8'h15;
mem[16'hBB1A] = 8'h7F;
mem[16'hBB1B] = 8'hBF;
mem[16'hBB1C] = 8'h20;
mem[16'hBB1D] = 8'hB2;
mem[16'hBB1E] = 8'hFE;
mem[16'hBB1F] = 8'h32;
mem[16'hBB20] = 8'h37;
mem[16'hBB21] = 8'h08;
mem[16'hBB22] = 8'h82;
mem[16'hBB23] = 8'h26;
mem[16'hBB24] = 8'h37;
mem[16'hBB25] = 8'hC1;
mem[16'hBB26] = 8'h23;
mem[16'hBB27] = 8'hD7;
mem[16'hBB28] = 8'hCC;
mem[16'hBB29] = 8'hA5;
mem[16'hBB2A] = 8'h67;
mem[16'hBB2B] = 8'h3B;
mem[16'hBB2C] = 8'hA0;
mem[16'hBB2D] = 8'h81;
mem[16'hBB2E] = 8'h37;
mem[16'hBB2F] = 8'h2E;
mem[16'hBB30] = 8'h94;
mem[16'hBB31] = 8'h3D;
mem[16'hBB32] = 8'h6E;
mem[16'hBB33] = 8'h9D;
mem[16'hBB34] = 8'hF8;
mem[16'hBB35] = 8'hB9;
mem[16'hBB36] = 8'h37;
mem[16'hBB37] = 8'h92;
mem[16'hBB38] = 8'h34;
mem[16'hBB39] = 8'h10;
mem[16'hBB3A] = 8'h9E;
mem[16'hBB3B] = 8'h32;
mem[16'hBB3C] = 8'h9C;
mem[16'hBB3D] = 8'h41;
mem[16'hBB3E] = 8'h9F;
mem[16'hBB3F] = 8'h3E;
mem[16'hBB40] = 8'hEF;
mem[16'hBB41] = 8'h4D;
mem[16'hBB42] = 8'h6B;
mem[16'hBB43] = 8'hEE;
mem[16'hBB44] = 8'h41;
mem[16'hBB45] = 8'hEB;
mem[16'hBB46] = 8'h6F;
mem[16'hBB47] = 8'hEC;
mem[16'hBB48] = 8'hA8;
mem[16'hBB49] = 8'hEA;
mem[16'hBB4A] = 8'h53;
mem[16'hBB4B] = 8'h62;
mem[16'hBB4C] = 8'h29;
mem[16'hBB4D] = 8'hE3;
mem[16'hBB4E] = 8'h52;
mem[16'hBB4F] = 8'hE4;
mem[16'hBB50] = 8'h6C;
mem[16'hBB51] = 8'hFC;
mem[16'hBB52] = 8'h57;
mem[16'hBB53] = 8'hB3;
mem[16'hBB54] = 8'h61;
mem[16'hBB55] = 8'h42;
mem[16'hBB56] = 8'h53;
mem[16'hBB57] = 8'h2B;
mem[16'hBB58] = 8'hF0;
mem[16'hBB59] = 8'hB9;
mem[16'hBB5A] = 8'h5E;
mem[16'hBB5B] = 8'h4C;
mem[16'hBB5C] = 8'h75;
mem[16'hBB5D] = 8'h38;
mem[16'hBB5E] = 8'hF6;
mem[16'hBB5F] = 8'h43;
mem[16'hBB60] = 8'hC8;
mem[16'hBB61] = 8'h81;
mem[16'hBB62] = 8'h79;
mem[16'hBB63] = 8'h74;
mem[16'hBB64] = 8'h0D;
mem[16'hBB65] = 8'h19;
mem[16'hBB66] = 8'hCE;
mem[16'hBB67] = 8'h87;
mem[16'hBB68] = 8'h14;
mem[16'hBB69] = 8'h7E;
mem[16'hBB6A] = 8'h57;
mem[16'hBB6B] = 8'h0E;
mem[16'hBB6C] = 8'hC6;
mem[16'hBB6D] = 8'h71;
mem[16'hBB6E] = 8'hC6;
mem[16'hBB6F] = 8'h8F;
mem[16'hBB70] = 8'hC3;
mem[16'hBB71] = 8'h60;
mem[16'hBB72] = 8'h1C;
mem[16'hBB73] = 8'h0F;
mem[16'hBB74] = 8'hDC;
mem[16'hBB75] = 8'h95;
mem[16'hBB76] = 8'hF5;
mem[16'hBB77] = 8'h66;
mem[16'hBB78] = 8'hE5;
mem[16'hBB79] = 8'h1C;
mem[16'hBB7A] = 8'hDE;
mem[16'hBB7B] = 8'h67;
mem[16'hBB7C] = 8'hD4;
mem[16'hBB7D] = 8'h9D;
mem[16'hBB7E] = 8'hED;
mem[16'hBB7F] = 8'h6E;
mem[16'hBB80] = 8'h85;
mem[16'hBB81] = 8'hFD;
mem[16'hBB82] = 8'h22;
mem[16'hBB83] = 8'h63;
mem[16'hBB84] = 8'h65;
mem[16'hBB85] = 8'h97;
mem[16'hBB86] = 8'hF8;
mem[16'hBB87] = 8'hEE;
mem[16'hBB88] = 8'hE6;
mem[16'hBB89] = 8'hEA;
mem[16'hBB8A] = 8'hE9;
mem[16'hBB8B] = 8'hF3;
mem[16'hBB8C] = 8'hE9;
mem[16'hBB8D] = 8'hEF;
mem[16'hBB8E] = 8'hE5;
mem[16'hBB8F] = 8'hEA;
mem[16'hBB90] = 8'h35;
mem[16'hBB91] = 8'hCD;
mem[16'hBB92] = 8'h3C;
mem[16'hBB93] = 8'h5F;
mem[16'hBB94] = 8'hBD;
mem[16'hBB95] = 8'h75;
mem[16'hBB96] = 8'h4A;
mem[16'hBB97] = 8'h84;
mem[16'hBB98] = 8'hF6;
mem[16'hBB99] = 8'h7C;
mem[16'hBB9A] = 8'h37;
mem[16'hBB9B] = 8'hB2;
mem[16'hBB9C] = 8'h36;
mem[16'hBB9D] = 8'h11;
mem[16'hBB9E] = 8'hB8;
mem[16'hBB9F] = 8'h8F;
mem[16'hBBA0] = 8'hA5;
mem[16'hBBA1] = 8'h09;
mem[16'hBBA2] = 8'h8B;
mem[16'hBBA3] = 8'h08;
mem[16'hBBA4] = 8'h44;
mem[16'hBBA5] = 8'hD1;
mem[16'hBBA6] = 8'hBC;
mem[16'hBBA7] = 8'hA2;
mem[16'hBBA8] = 8'h4D;
mem[16'hBBA9] = 8'h07;
mem[16'hBBAA] = 8'h83;
mem[16'hBBAB] = 8'h01;
mem[16'hBBAC] = 8'h20;
mem[16'hBBAD] = 8'h8B;
mem[16'hBBAE] = 8'hBE;
mem[16'hBBAF] = 8'hAA;
mem[16'hBBB0] = 8'h1A;
mem[16'hBBB1] = 8'h98;
mem[16'hBBB2] = 8'h19;
mem[16'hBBB3] = 8'h53;
mem[16'hBBB4] = 8'h18;
mem[16'hBBB5] = 8'hA0;
mem[16'hBBB6] = 8'h9F;
mem[16'hBBB7] = 8'h52;
mem[16'hBBB8] = 8'h17;
mem[16'hBBB9] = 8'h90;
mem[16'hBBBA] = 8'h10;
mem[16'hBBBB] = 8'h37;
mem[16'hBBBC] = 8'h9A;
mem[16'hBBBD] = 8'hAD;
mem[16'hBBBE] = 8'hBB;
mem[16'hBBBF] = 8'hBB;
mem[16'hBBC0] = 8'hCC;
mem[16'hBBC1] = 8'h6D;
mem[16'hBBC2] = 8'hF7;
mem[16'hBBC3] = 8'h6F;
mem[16'hBBC4] = 8'hC1;
mem[16'hBBC5] = 8'hA1;
mem[16'hBBC6] = 8'hBA;
mem[16'hBBC7] = 8'h91;
mem[16'hBBC8] = 8'hCD;
mem[16'hBBC9] = 8'h61;
mem[16'hBBCA] = 8'hE3;
mem[16'hBBCB] = 8'h60;
mem[16'hBBCC] = 8'h2C;
mem[16'hBBCD] = 8'hB9;
mem[16'hBBCE] = 8'hD4;
mem[16'hBBCF] = 8'hCA;
mem[16'hBBD0] = 8'h35;
mem[16'hBBD1] = 8'h79;
mem[16'hBBD2] = 8'hFB;
mem[16'hBBD3] = 8'h79;
mem[16'hBBD4] = 8'hD5;
mem[16'hBBD5] = 8'h73;
mem[16'hBBD6] = 8'hDA;
mem[16'hBBD7] = 8'hFE;
mem[16'hBBD8] = 8'h7F;
mem[16'hBBD9] = 8'hD5;
mem[16'hBBDA] = 8'h76;
mem[16'hBBDB] = 8'hEF;
mem[16'hBBDC] = 8'hE9;
mem[16'hBBDD] = 8'h71;
mem[16'hBBDE] = 8'hDA;
mem[16'hBBDF] = 8'hBB;
mem[16'hBBE0] = 8'h9C;
mem[16'hBBE1] = 8'hB7;
mem[16'hBBE2] = 8'hE7;
mem[16'hBBE3] = 8'hD7;
mem[16'hBBE4] = 8'hCD;
mem[16'hBBE5] = 8'h49;
mem[16'hBBE6] = 8'hE3;
mem[16'hBBE7] = 8'h4B;
mem[16'hBBE8] = 8'hC1;
mem[16'hBBE9] = 8'h44;
mem[16'hBBEA] = 8'h66;
mem[16'hBBEB] = 8'h48;
mem[16'hBBEC] = 8'hF5;
mem[16'hBBED] = 8'hEC;
mem[16'hBBEE] = 8'h47;
mem[16'hBBEF] = 8'hE3;
mem[16'hBBF0] = 8'hAC;
mem[16'hBBF1] = 8'h56;
mem[16'hBBF2] = 8'h97;
mem[16'hBBF3] = 8'h5B;
mem[16'hBBF4] = 8'hE8;
mem[16'hBBF5] = 8'h55;
mem[16'hBBF6] = 8'hF3;
mem[16'hBBF7] = 8'h5E;
mem[16'hBBF8] = 8'hD9;
mem[16'hBBF9] = 8'h5D;
mem[16'hBBFA] = 8'hF6;
mem[16'hBBFB] = 8'h37;
mem[16'hBBFC] = 8'hD5;
mem[16'hBBFD] = 8'hF8;
mem[16'hBBFE] = 8'h56;
mem[16'hBBFF] = 8'hDE;
mem[16'hBC00] = 8'hA9;
mem[16'hBC01] = 8'h0D;
mem[16'hBC02] = 8'h0E;
mem[16'hBC03] = 8'hAF;
mem[16'hBC04] = 8'h05;
mem[16'hBC05] = 8'hAA;
mem[16'hBC06] = 8'h0A;
mem[16'hBC07] = 8'h2E;
mem[16'hBC08] = 8'hA5;
mem[16'hBC09] = 8'h85;
mem[16'hBC0A] = 8'hEA;
mem[16'hBC0B] = 8'h1B;
mem[16'hBC0C] = 8'h66;
mem[16'hBC0D] = 8'hAA;
mem[16'hBC0E] = 8'h52;
mem[16'hBC0F] = 8'hB3;
mem[16'hBC10] = 8'h19;
mem[16'hBC11] = 8'hBC;
mem[16'hBC12] = 8'hA6;
mem[16'hBC13] = 8'hD2;
mem[16'hBC14] = 8'hBD;
mem[16'hBC15] = 8'h19;
mem[16'hBC16] = 8'h2A;
mem[16'hBC17] = 8'hB9;
mem[16'hBC18] = 8'h1D;
mem[16'hBC19] = 8'h4A;
mem[16'hBC1A] = 8'h33;
mem[16'hBC1B] = 8'hB6;
mem[16'hBC1C] = 8'h79;
mem[16'hBC1D] = 8'h3D;
mem[16'hBC1E] = 8'h02;
mem[16'hBC1F] = 8'hB3;
mem[16'hBC20] = 8'h25;
mem[16'hBC21] = 8'h9D;
mem[16'hBC22] = 8'h0B;
mem[16'hBC23] = 8'h94;
mem[16'hBC24] = 8'h21;
mem[16'hBC25] = 8'h8F;
mem[16'hBC26] = 8'h0F;
mem[16'hBC27] = 8'h8C;
mem[16'hBC28] = 8'h21;
mem[16'hBC29] = 8'h84;
mem[16'hBC2A] = 8'hCE;
mem[16'hBC2B] = 8'hA7;
mem[16'hBC2C] = 8'h83;
mem[16'hBC2D] = 8'h38;
mem[16'hBC2E] = 8'hEA;
mem[16'hBC2F] = 8'h06;
mem[16'hBC30] = 8'h9D;
mem[16'hBC31] = 8'h34;
mem[16'hBC32] = 8'hC8;
mem[16'hBC33] = 8'h1A;
mem[16'hBC34] = 8'h83;
mem[16'hBC35] = 8'h34;
mem[16'hBC36] = 8'h92;
mem[16'hBC37] = 8'h3B;
mem[16'hBC38] = 8'h64;
mem[16'hBC39] = 8'h97;
mem[16'hBC3A] = 8'hF6;
mem[16'hBC3B] = 8'hB7;
mem[16'hBC3C] = 8'h35;
mem[16'hBC3D] = 8'h90;
mem[16'hBC3E] = 8'h5B;
mem[16'hBC3F] = 8'h1F;
mem[16'hBC40] = 8'h5C;
mem[16'hBC41] = 8'hE5;
mem[16'hBC42] = 8'h4E;
mem[16'hBC43] = 8'hEF;
mem[16'hBC44] = 8'h4D;
mem[16'hBC45] = 8'hE2;
mem[16'hBC46] = 8'h3A;
mem[16'hBC47] = 8'h2A;
mem[16'hBC48] = 8'h84;
mem[16'hBC49] = 8'hB0;
mem[16'hBC4A] = 8'h86;
mem[16'hBC4B] = 8'hC7;
mem[16'hBC4C] = 8'h78;
mem[16'hBC4D] = 8'hC8;
mem[16'hBC4E] = 8'hED;
mem[16'hBC4F] = 8'h66;
mem[16'hBC50] = 8'hF9;
mem[16'hBC51] = 8'h54;
mem[16'hBC52] = 8'h56;
mem[16'hBC53] = 8'h7A;
mem[16'hBC54] = 8'hF0;
mem[16'hBC55] = 8'hD9;
mem[16'hBC56] = 8'h9A;
mem[16'hBC57] = 8'h47;
mem[16'hBC58] = 8'h3C;
mem[16'hBC59] = 8'h6D;
mem[16'hBC5A] = 8'hDF;
mem[16'hBC5B] = 8'hF8;
mem[16'hBC5C] = 8'h20;
mem[16'hBC5D] = 8'h00;
mem[16'hBC5E] = 8'h92;
mem[16'hBC5F] = 8'h5A;
mem[16'hBC60] = 8'h69;
mem[16'hBC61] = 8'hC8;
mem[16'hBC62] = 8'hC4;
mem[16'hBC63] = 8'hC5;
mem[16'hBC64] = 8'h8D;
mem[16'hBC65] = 8'hC8;
mem[16'hBC66] = 8'hE3;
mem[16'hBC67] = 8'hF4;
mem[16'hBC68] = 8'h6E;
mem[16'hBC69] = 8'h78;
mem[16'hBC6A] = 8'hC6;
mem[16'hBC6B] = 8'h6B;
mem[16'hBC6C] = 8'h59;
mem[16'hBC6D] = 8'hC1;
mem[16'hBC6E] = 8'h69;
mem[16'hBC6F] = 8'h66;
mem[16'hBC70] = 8'hD4;
mem[16'hBC71] = 8'h44;
mem[16'hBC72] = 8'hDE;
mem[16'hBC73] = 8'h76;
mem[16'hBC74] = 8'h7D;
mem[16'hBC75] = 8'hD8;
mem[16'hBC76] = 8'h43;
mem[16'hBC77] = 8'hDB;
mem[16'hBC78] = 8'h7E;
mem[16'hBC79] = 8'h1D;
mem[16'hBC7A] = 8'h26;
mem[16'hBC7B] = 8'hDC;
mem[16'hBC7C] = 8'h79;
mem[16'hBC7D] = 8'h2E;
mem[16'hBC7E] = 8'h4B;
mem[16'hBC7F] = 8'hD3;
mem[16'hBC80] = 8'h85;
mem[16'hBC81] = 8'hB4;
mem[16'hBC82] = 8'h2E;
mem[16'hBC83] = 8'h85;
mem[16'hBC84] = 8'hB1;
mem[16'hBC85] = 8'h29;
mem[16'hBC86] = 8'h81;
mem[16'hBC87] = 8'hA3;
mem[16'hBC88] = 8'h44;
mem[16'hBC89] = 8'hB0;
mem[16'hBC8A] = 8'h8B;
mem[16'hBC8B] = 8'h23;
mem[16'hBC8C] = 8'h80;
mem[16'hBC8D] = 8'hA4;
mem[16'hBC8E] = 8'h27;
mem[16'hBC8F] = 8'h8E;
mem[16'hBC90] = 8'h39;
mem[16'hBC91] = 8'h9D;
mem[16'hBC92] = 8'hEE;
mem[16'hBC93] = 8'h37;
mem[16'hBC94] = 8'h91;
mem[16'hBC95] = 8'h3D;
mem[16'hBC96] = 8'hB7;
mem[16'hBC97] = 8'h3E;
mem[16'hBC98] = 8'h94;
mem[16'hBC99] = 8'h79;
mem[16'hBC9A] = 8'h9E;
mem[16'hBC9B] = 8'h8B;
mem[16'hBC9C] = 8'hF9;
mem[16'hBC9D] = 8'h35;
mem[16'hBC9E] = 8'h82;
mem[16'hBC9F] = 8'h3B;
mem[16'hBCA0] = 8'hA5;
mem[16'hBCA1] = 8'h08;
mem[16'hBCA2] = 8'h83;
mem[16'hBCA3] = 8'h07;
mem[16'hBCA4] = 8'hA8;
mem[16'hBCA5] = 8'h61;
mem[16'hBCA6] = 8'h62;
mem[16'hBCA7] = 8'h6B;
mem[16'hBCA8] = 8'hA9;
mem[16'hBCA9] = 8'h0F;
mem[16'hBCAA] = 8'hA6;
mem[16'hBCAB] = 8'h82;
mem[16'hBCAC] = 8'h0F;
mem[16'hBCAD] = 8'hAC;
mem[16'hBCAE] = 8'h0B;
mem[16'hBCAF] = 8'hA3;
mem[16'hBCB0] = 8'h99;
mem[16'hBCB1] = 8'h15;
mem[16'hBCB2] = 8'hB3;
mem[16'hBCB3] = 8'h1C;
mem[16'hBCB4] = 8'hB8;
mem[16'hBCB5] = 8'h9C;
mem[16'hBCB6] = 8'h1B;
mem[16'hBCB7] = 8'hBB;
mem[16'hBCB8] = 8'h14;
mem[16'hBCB9] = 8'h35;
mem[16'hBCBA] = 8'h76;
mem[16'hBCBB] = 8'hAB;
mem[16'hBCBC] = 8'hD6;
mem[16'hBCBD] = 8'h1E;
mem[16'hBCBE] = 8'hE2;
mem[16'hBCBF] = 8'h33;
mem[16'hBCC0] = 8'hA4;
mem[16'hBCC1] = 8'h8B;
mem[16'hBCC2] = 8'h66;
mem[16'hBCC3] = 8'h89;
mem[16'hBCC4] = 8'h6D;
mem[16'hBCC5] = 8'hCC;
mem[16'hBCC6] = 8'h6F;
mem[16'hBCC7] = 8'h42;
mem[16'hBCC8] = 8'h6B;
mem[16'hBCC9] = 8'hB5;
mem[16'hBCCA] = 8'h88;
mem[16'hBCCB] = 8'hE2;
mem[16'hBCCC] = 8'h65;
mem[16'hBCCD] = 8'hC4;
mem[16'hBCCE] = 8'h63;
mem[16'hBCCF] = 8'h7B;
mem[16'hBCD0] = 8'h11;
mem[16'hBCD1] = 8'h78;
mem[16'hBCD2] = 8'hDE;
mem[16'hBCD3] = 8'hFA;
mem[16'hBCD4] = 8'h79;
mem[16'hBCD5] = 8'hB0;
mem[16'hBCD6] = 8'hF6;
mem[16'hBCD7] = 8'hEB;
mem[16'hBCD8] = 8'h94;
mem[16'hBCD9] = 8'hDC;
mem[16'hBCDA] = 8'h7C;
mem[16'hBCDB] = 8'hFA;
mem[16'hBCDC] = 8'h78;
mem[16'hBCDD] = 8'hD1;
mem[16'hBCDE] = 8'h1A;
mem[16'hBCDF] = 8'h1B;
mem[16'hBCE0] = 8'h2C;
mem[16'hBCE1] = 8'hE0;
mem[16'hBCE2] = 8'h4F;
mem[16'hBCE3] = 8'hEF;
mem[16'hBCE4] = 8'h61;
mem[16'hBCE5] = 8'h39;
mem[16'hBCE6] = 8'h9A;
mem[16'hBCE7] = 8'h42;
mem[16'hBCE8] = 8'hED;
mem[16'hBCE9] = 8'h44;
mem[16'hBCEA] = 8'hCB;
mem[16'hBCEB] = 8'h4F;
mem[16'hBCEC] = 8'hE0;
mem[16'hBCED] = 8'h29;
mem[16'hBCEE] = 8'h2A;
mem[16'hBCEF] = 8'h23;
mem[16'hBCF0] = 8'hF5;
mem[16'hBCF1] = 8'hD8;
mem[16'hBCF2] = 8'h54;
mem[16'hBCF3] = 8'h15;
mem[16'hBCF4] = 8'h12;
mem[16'hBCF5] = 8'h13;
mem[16'hBCF6] = 8'hF2;
mem[16'hBCF7] = 8'hF6;
mem[16'hBCF8] = 8'h56;
mem[16'hBCF9] = 8'hF5;
mem[16'hBCFA] = 8'hA6;
mem[16'hBCFB] = 8'h53;
mem[16'hBCFC] = 8'h99;
mem[16'hBCFD] = 8'h52;
mem[16'hBCFE] = 8'hC2;
mem[16'hBCFF] = 8'h5B;
mem[16'hBD00] = 8'h05;
mem[16'hBD01] = 8'hAF;
mem[16'hBD02] = 8'h23;
mem[16'hBD03] = 8'hA7;
mem[16'hBD04] = 8'h08;
mem[16'hBD05] = 8'hC1;
mem[16'hBD06] = 8'hC2;
mem[16'hBD07] = 8'hCB;
mem[16'hBD08] = 8'h21;
mem[16'hBD09] = 8'hAE;
mem[16'hBD0A] = 8'h6F;
mem[16'hBD0B] = 8'hA5;
mem[16'hBD0C] = 8'h30;
mem[16'hBD0D] = 8'hA0;
mem[16'hBD0E] = 8'h6A;
mem[16'hBD0F] = 8'h1A;
mem[16'hBD10] = 8'h4C;
mem[16'hBD11] = 8'h09;
mem[16'hBD12] = 8'h3B;
mem[16'hBD13] = 8'hBF;
mem[16'hBD14] = 8'h35;
mem[16'hBD15] = 8'hB9;
mem[16'hBD16] = 8'h1A;
mem[16'hBD17] = 8'h3F;
mem[16'hBD18] = 8'hAD;
mem[16'hBD19] = 8'h1C;
mem[16'hBD1A] = 8'hE0;
mem[16'hBD1B] = 8'h32;
mem[16'hBD1C] = 8'hAB;
mem[16'hBD1D] = 8'hD1;
mem[16'hBD1E] = 8'h9B;
mem[16'hBD1F] = 8'h1A;
mem[16'hBD20] = 8'h3A;
mem[16'hBD21] = 8'h08;
mem[16'hBD22] = 8'h9B;
mem[16'hBD23] = 8'h26;
mem[16'hBD24] = 8'h50;
mem[16'hBD25] = 8'h0C;
mem[16'hBD26] = 8'h9E;
mem[16'hBD27] = 8'h22;
mem[16'hBD28] = 8'h84;
mem[16'hBD29] = 8'h00;
mem[16'hBD2A] = 8'h81;
mem[16'hBD2B] = 8'hCB;
mem[16'hBD2C] = 8'hE2;
mem[16'hBD2D] = 8'h3C;
mem[16'hBD2E] = 8'hCB;
mem[16'hBD2F] = 8'h2A;
mem[16'hBD30] = 8'h25;
mem[16'hBD31] = 8'h18;
mem[16'hBD32] = 8'h8B;
mem[16'hBD33] = 8'h36;
mem[16'hBD34] = 8'h98;
mem[16'hBD35] = 8'h1C;
mem[16'hBD36] = 8'h8E;
mem[16'hBD37] = 8'h32;
mem[16'hBD38] = 8'h92;
mem[16'hBD39] = 8'h10;
mem[16'hBD3A] = 8'h91;
mem[16'hBD3B] = 8'hDB;
mem[16'hBD3C] = 8'hF2;
mem[16'hBD3D] = 8'h2C;
mem[16'hBD3E] = 8'h8B;
mem[16'hBD3F] = 8'h3A;
mem[16'hBD40] = 8'h51;
mem[16'hBD41] = 8'h68;
mem[16'hBD42] = 8'hFB;
mem[16'hBD43] = 8'h46;
mem[16'hBD44] = 8'hA7;
mem[16'hBD45] = 8'h6C;
mem[16'hBD46] = 8'hFE;
mem[16'hBD47] = 8'h42;
mem[16'hBD48] = 8'hE4;
mem[16'hBD49] = 8'h60;
mem[16'hBD4A] = 8'hE1;
mem[16'hBD4B] = 8'hAB;
mem[16'hBD4C] = 8'h82;
mem[16'hBD4D] = 8'h5C;
mem[16'hBD4E] = 8'h8B;
mem[16'hBD4F] = 8'h41;
mem[16'hBD50] = 8'hFC;
mem[16'hBD51] = 8'h40;
mem[16'hBD52] = 8'hFE;
mem[16'hBD53] = 8'h56;
mem[16'hBD54] = 8'h08;
mem[16'hBD55] = 8'hFC;
mem[16'hBD56] = 8'h53;
mem[16'hBD57] = 8'h53;
mem[16'hBD58] = 8'h69;
mem[16'hBD59] = 8'hF5;
mem[16'hBD5A] = 8'h5F;
mem[16'hBD5B] = 8'h1F;
mem[16'hBD5C] = 8'h20;
mem[16'hBD5D] = 8'h02;
mem[16'hBD5E] = 8'hBE;
mem[16'hBD5F] = 8'h2B;
mem[16'hBD60] = 8'h7A;
mem[16'hBD61] = 8'hB4;
mem[16'hBD62] = 8'h60;
mem[16'hBD63] = 8'hC9;
mem[16'hBD64] = 8'h68;
mem[16'hBD65] = 8'h29;
mem[16'hBD66] = 8'hDA;
mem[16'hBD67] = 8'h5B;
mem[16'hBD68] = 8'hC2;
mem[16'hBD69] = 8'h6C;
mem[16'hBD6A] = 8'hC0;
mem[16'hBD6B] = 8'h4A;
mem[16'hBD6C] = 8'hC8;
mem[16'hBD6D] = 8'h61;
mem[16'hBD6E] = 8'hA2;
mem[16'hBD6F] = 8'h6E;
mem[16'hBD70] = 8'hD5;
mem[16'hBD71] = 8'h7D;
mem[16'hBD72] = 8'h0E;
mem[16'hBD73] = 8'hDC;
mem[16'hBD74] = 8'h65;
mem[16'hBD75] = 8'hD9;
mem[16'hBD76] = 8'h68;
mem[16'hBD77] = 8'h5E;
mem[16'hBD78] = 8'hDC;
mem[16'hBD79] = 8'h7C;
mem[16'hBD7A] = 8'hD6;
mem[16'hBD7B] = 8'h52;
mem[16'hBD7C] = 8'hD9;
mem[16'hBD7D] = 8'hF1;
mem[16'hBD7E] = 8'h4B;
mem[16'hBD7F] = 8'h6E;
mem[16'hBD80] = 8'h0C;
mem[16'hBD81] = 8'hC7;
mem[16'hBD82] = 8'h93;
mem[16'hBD83] = 8'h82;
mem[16'hBD84] = 8'h20;
mem[16'hBD85] = 8'h89;
mem[16'hBD86] = 8'hFA;
mem[16'hBD87] = 8'h20;
mem[16'hBD88] = 8'h81;
mem[16'hBD89] = 8'h2C;
mem[16'hBD8A] = 8'h3E;
mem[16'hBD8B] = 8'h4E;
mem[16'hBD8C] = 8'h10;
mem[16'hBD8D] = 8'hA4;
mem[16'hBD8E] = 8'h2B;
mem[16'hBD8F] = 8'hEA;
mem[16'hBD90] = 8'hFC;
mem[16'hBD91] = 8'hAD;
mem[16'hBD92] = 8'hD4;
mem[16'hBD93] = 8'h5F;
mem[16'hBD94] = 8'h74;
mem[16'hBD95] = 8'h55;
mem[16'hBD96] = 8'h2E;
mem[16'hBD97] = 8'h3B;
mem[16'hBD98] = 8'h3D;
mem[16'hBD99] = 8'h95;
mem[16'hBD9A] = 8'hBD;
mem[16'hBD9B] = 8'h9E;
mem[16'hBD9C] = 8'hB1;
mem[16'hBD9D] = 8'hA8;
mem[16'hBD9E] = 8'h32;
mem[16'hBD9F] = 8'h9B;
mem[16'hBDA0] = 8'h84;
mem[16'hBDA1] = 8'hDD;
mem[16'hBDA2] = 8'hF4;
mem[16'hBDA3] = 8'h82;
mem[16'hBDA4] = 8'h08;
mem[16'hBDA5] = 8'hA1;
mem[16'hBDA6] = 8'hA8;
mem[16'hBDA7] = 8'h04;
mem[16'hBDA8] = 8'hB9;
mem[16'hBDA9] = 8'h85;
mem[16'hBDAA] = 8'hB5;
mem[16'hBDAB] = 8'hF7;
mem[16'hBDAC] = 8'h38;
mem[16'hBDAD] = 8'hC8;
mem[16'hBDAE] = 8'h01;
mem[16'hBDAF] = 8'hB3;
mem[16'hBDB0] = 8'h28;
mem[16'hBDB1] = 8'h17;
mem[16'hBDB2] = 8'hD7;
mem[16'hBDB3] = 8'h1D;
mem[16'hBDB4] = 8'hE8;
mem[16'hBDB5] = 8'h18;
mem[16'hBDB6] = 8'h10;
mem[16'hBDB7] = 8'h9E;
mem[16'hBDB8] = 8'h04;
mem[16'hBDB9] = 8'h9F;
mem[16'hBDBA] = 8'h1C;
mem[16'hBDBB] = 8'h1D;
mem[16'hBDBC] = 8'h1A;
mem[16'hBDBD] = 8'h1B;
mem[16'hBDBE] = 8'h17;
mem[16'hBDBF] = 8'h03;
mem[16'hBDC0] = 8'hE9;
mem[16'hBDC1] = 8'h7D;
mem[16'hBDC2] = 8'hD2;
mem[16'hBDC3] = 8'hFF;
mem[16'hBDC4] = 8'hDB;
mem[16'hBDC5] = 8'hCC;
mem[16'hBDC6] = 8'h7A;
mem[16'hBDC7] = 8'hF2;
mem[16'hBDC8] = 8'h64;
mem[16'hBDC9] = 8'hCD;
mem[16'hBDCA] = 8'hC3;
mem[16'hBDCB] = 8'h77;
mem[16'hBDCC] = 8'h49;
mem[16'hBDCD] = 8'h69;
mem[16'hBDCE] = 8'hB2;
mem[16'hBDCF] = 8'h60;
mem[16'hBDD0] = 8'hB4;
mem[16'hBDD1] = 8'hAD;
mem[16'hBDD2] = 8'h74;
mem[16'hBDD3] = 8'hE7;
mem[16'hBDD4] = 8'h60;
mem[16'hBDD5] = 8'h04;
mem[16'hBDD6] = 8'hCA;
mem[16'hBDD7] = 8'hC8;
mem[16'hBDD8] = 8'hDC;
mem[16'hBDD9] = 8'hE5;
mem[16'hBDDA] = 8'h74;
mem[16'hBDDB] = 8'hD7;
mem[16'hBDDC] = 8'h8F;
mem[16'hBDDD] = 8'hE9;
mem[16'hBDDE] = 8'hAF;
mem[16'hBDDF] = 8'hD3;
mem[16'hBDE0] = 8'hFF;
mem[16'hBDE1] = 8'hDD;
mem[16'hBDE2] = 8'hAC;
mem[16'hBDE3] = 8'hBF;
mem[16'hBDE4] = 8'hA8;
mem[16'hBDE5] = 8'h83;
mem[16'hBDE6] = 8'h5A;
mem[16'hBDE7] = 8'h8B;
mem[16'hBDE8] = 8'h24;
mem[16'hBDE9] = 8'hBC;
mem[16'hBDEA] = 8'hE3;
mem[16'hBDEB] = 8'h4E;
mem[16'hBDEC] = 8'h58;
mem[16'hBDED] = 8'h4C;
mem[16'hBDEE] = 8'h44;
mem[16'hBDEF] = 8'hE3;
mem[16'hBDF0] = 8'hF6;
mem[16'hBDF1] = 8'hE0;
mem[16'hBDF2] = 8'h1E;
mem[16'hBDF3] = 8'hED;
mem[16'hBDF4] = 8'h88;
mem[16'hBDF5] = 8'h58;
mem[16'hBDF6] = 8'h3A;
mem[16'hBDF7] = 8'hDE;
mem[16'hBDF8] = 8'h45;
mem[16'hBDF9] = 8'hC5;
mem[16'hBDFA] = 8'h54;
mem[16'hBDFB] = 8'h37;
mem[16'hBDFC] = 8'h1C;
mem[16'hBDFD] = 8'hEC;
mem[16'hBDFE] = 8'h62;
mem[16'hBDFF] = 8'hE1;
mem[16'hBE00] = 8'h29;
mem[16'hBE01] = 8'hA8;
mem[16'hBE02] = 8'h0E;
mem[16'hBE03] = 8'hAF;
mem[16'hBE04] = 8'h15;
mem[16'hBE05] = 8'h89;
mem[16'hBE06] = 8'h18;
mem[16'hBE07] = 8'h01;
mem[16'hBE08] = 8'h22;
mem[16'hBE09] = 8'hA4;
mem[16'hBE0A] = 8'h86;
mem[16'hBE0B] = 8'hC7;
mem[16'hBE0C] = 8'h1C;
mem[16'hBE0D] = 8'h47;
mem[16'hBE0E] = 8'hAA;
mem[16'hBE0F] = 8'h65;
mem[16'hBE10] = 8'hAD;
mem[16'hBE11] = 8'h4D;
mem[16'hBE12] = 8'h88;
mem[16'hBE13] = 8'h77;
mem[16'hBE14] = 8'h5E;
mem[16'hBE15] = 8'hBC;
mem[16'hBE16] = 8'h1C;
mem[16'hBE17] = 8'hBA;
mem[16'hBE18] = 8'h09;
mem[16'hBE19] = 8'hB5;
mem[16'hBE1A] = 8'h1E;
mem[16'hBE1B] = 8'h9E;
mem[16'hBE1C] = 8'hBF;
mem[16'hBE1D] = 8'hBB;
mem[16'hBE1E] = 8'h37;
mem[16'hBE1F] = 8'hA3;
mem[16'hBE20] = 8'h29;
mem[16'hBE21] = 8'h88;
mem[16'hBE22] = 8'h4B;
mem[16'hBE23] = 8'h9F;
mem[16'hBE24] = 8'h18;
mem[16'hBE25] = 8'h6D;
mem[16'hBE26] = 8'h23;
mem[16'hBE27] = 8'h8B;
mem[16'hBE28] = 8'h01;
mem[16'hBE29] = 8'h80;
mem[16'hBE2A] = 8'h23;
mem[16'hBE2B] = 8'h97;
mem[16'hBE2C] = 8'h49;
mem[16'hBE2D] = 8'h91;
mem[16'hBE2E] = 8'h32;
mem[16'hBE2F] = 8'h86;
mem[16'hBE30] = 8'h74;
mem[16'hBE31] = 8'h1B;
mem[16'hBE32] = 8'h9F;
mem[16'hBE33] = 8'h4F;
mem[16'hBE34] = 8'h4D;
mem[16'hBE35] = 8'h24;
mem[16'hBE36] = 8'h9A;
mem[16'hBE37] = 8'h33;
mem[16'hBE38] = 8'hDE;
mem[16'hBE39] = 8'hDF;
mem[16'hBE3A] = 8'hDC;
mem[16'hBE3B] = 8'hDD;
mem[16'hBE3C] = 8'h3A;
mem[16'hBE3D] = 8'h2C;
mem[16'hBE3E] = 8'h22;
mem[16'hBE3F] = 8'h20;
mem[16'hBE40] = 8'hF4;
mem[16'hBE41] = 8'h88;
mem[16'hBE42] = 8'hEF;
mem[16'hBE43] = 8'h6A;
mem[16'hBE44] = 8'hE9;
mem[16'hBE45] = 8'h43;
mem[16'hBE46] = 8'h3A;
mem[16'hBE47] = 8'h29;
mem[16'hBE48] = 8'hC4;
mem[16'hBE49] = 8'hA9;
mem[16'hBE4A] = 8'h73;
mem[16'hBE4B] = 8'h5A;
mem[16'hBE4C] = 8'h69;
mem[16'hBE4D] = 8'h43;
mem[16'hBE4E] = 8'hE5;
mem[16'hBE4F] = 8'h69;
mem[16'hBE50] = 8'hF5;
mem[16'hBE51] = 8'h3D;
mem[16'hBE52] = 8'h7B;
mem[16'hBE53] = 8'hEE;
mem[16'hBE54] = 8'h58;
mem[16'hBE55] = 8'hF9;
mem[16'hBE56] = 8'h7E;
mem[16'hBE57] = 8'hEB;
mem[16'hBE58] = 8'h54;
mem[16'hBE59] = 8'hE5;
mem[16'hBE5A] = 8'h5F;
mem[16'hBE5B] = 8'hF0;
mem[16'hBE5C] = 8'h75;
mem[16'hBE5D] = 8'hFC;
mem[16'hBE5E] = 8'h43;
mem[16'hBE5F] = 8'hE3;
mem[16'hBE60] = 8'h49;
mem[16'hBE61] = 8'hC6;
mem[16'hBE62] = 8'h82;
mem[16'hBE63] = 8'hA8;
mem[16'hBE64] = 8'h76;
mem[16'hBE65] = 8'h78;
mem[16'hBE66] = 8'hDA;
mem[16'hBE67] = 8'h1A;
mem[16'hBE68] = 8'hD4;
mem[16'hBE69] = 8'h15;
mem[16'hBE6A] = 8'hD7;
mem[16'hBE6B] = 8'h16;
mem[16'hBE6C] = 8'hD0;
mem[16'hBE6D] = 8'h11;
mem[16'hBE6E] = 8'hCF;
mem[16'hBE6F] = 8'h06;
mem[16'hBE70] = 8'hD7;
mem[16'hBE71] = 8'h0D;
mem[16'hBE72] = 8'hDA;
mem[16'hBE73] = 8'h19;
mem[16'hBE74] = 8'hD5;
mem[16'hBE75] = 8'h29;
mem[16'hBE76] = 8'hDF;
mem[16'hBE77] = 8'h53;
mem[16'hBE78] = 8'hC4;
mem[16'hBE79] = 8'h3E;
mem[16'hBE7A] = 8'hE6;
mem[16'hBE7B] = 8'hD2;
mem[16'hBE7C] = 8'h79;
mem[16'hBE7D] = 8'hD1;
mem[16'hBE7E] = 8'h7A;
mem[16'hBE7F] = 8'h23;
mem[16'hBE80] = 8'h24;
mem[16'hBE81] = 8'h8D;
mem[16'hBE82] = 8'h2E;
mem[16'hBE83] = 8'hB7;
mem[16'hBE84] = 8'h79;
mem[16'hBE85] = 8'h39;
mem[16'hBE86] = 8'hE2;
mem[16'hBE87] = 8'hFB;
mem[16'hBE88] = 8'hDF;
mem[16'hBE89] = 8'hB8;
mem[16'hBE8A] = 8'h36;
mem[16'hBE8B] = 8'h87;
mem[16'hBE8C] = 8'hFD;
mem[16'hBE8D] = 8'hC1;
mem[16'hBE8E] = 8'h96;
mem[16'hBE8F] = 8'hD3;
mem[16'hBE90] = 8'h3F;
mem[16'hBE91] = 8'hD3;
mem[16'hBE92] = 8'h36;
mem[16'hBE93] = 8'h9F;
mem[16'hBE94] = 8'hF2;
mem[16'hBE95] = 8'hE9;
mem[16'hBE96] = 8'h82;
mem[16'hBE97] = 8'h96;
mem[16'hBE98] = 8'hB7;
mem[16'hBE99] = 8'hF5;
mem[16'hBE9A] = 8'h9B;
mem[16'hBE9B] = 8'hB4;
mem[16'hBE9C] = 8'hF0;
mem[16'hBE9D] = 8'h9C;
mem[16'hBE9E] = 8'h32;
mem[16'hBE9F] = 8'hD3;
mem[16'hBEA0] = 8'hAC;
mem[16'hBEA1] = 8'hF2;
mem[16'hBEA2] = 8'h82;
mem[16'hBEA3] = 8'h0F;
mem[16'hBEA4] = 8'hE8;
mem[16'hBEA5] = 8'hC5;
mem[16'hBEA6] = 8'h0A;
mem[16'hBEA7] = 8'hEB;
mem[16'hBEA8] = 8'hD4;
mem[16'hBEA9] = 8'h07;
mem[16'hBEAA] = 8'hC0;
mem[16'hBEAB] = 8'h17;
mem[16'hBEAC] = 8'h8D;
mem[16'hBEAD] = 8'h01;
mem[16'hBEAE] = 8'hE2;
mem[16'hBEAF] = 8'hAE;
mem[16'hBEB0] = 8'h9C;
mem[16'hBEB1] = 8'hDD;
mem[16'hBEB2] = 8'hBB;
mem[16'hBEB3] = 8'h0F;
mem[16'hBEB4] = 8'h31;
mem[16'hBEB5] = 8'h3B;
mem[16'hBEB6] = 8'h9F;
mem[16'hBEB7] = 8'h16;
mem[16'hBEB8] = 8'hC4;
mem[16'hBEB9] = 8'h22;
mem[16'hBEBA] = 8'hBF;
mem[16'hBEBB] = 8'hEF;
mem[16'hBEBC] = 8'h30;
mem[16'hBEBD] = 8'h57;
mem[16'hBEBE] = 8'hAD;
mem[16'hBEBF] = 8'hDA;
mem[16'hBEC0] = 8'hD5;
mem[16'hBEC1] = 8'hBD;
mem[16'hBEC2] = 8'h66;
mem[16'hBEC3] = 8'hCA;
mem[16'hBEC4] = 8'h65;
mem[16'hBEC5] = 8'h60;
mem[16'hBEC6] = 8'h6B;
mem[16'hBEC7] = 8'hEE;
mem[16'hBEC8] = 8'h69;
mem[16'hBEC9] = 8'hB5;
mem[16'hBECA] = 8'h6C;
mem[16'hBECB] = 8'hAE;
mem[16'hBECC] = 8'hF6;
mem[16'hBECD] = 8'h91;
mem[16'hBECE] = 8'h64;
mem[16'hBECF] = 8'hC6;
mem[16'hBED0] = 8'h71;
mem[16'hBED1] = 8'h74;
mem[16'hBED2] = 8'h7D;
mem[16'hBED3] = 8'hFA;
mem[16'hBED4] = 8'h75;
mem[16'hBED5] = 8'hD4;
mem[16'hBED6] = 8'hFA;
mem[16'hBED7] = 8'hBB;
mem[16'hBED8] = 8'hDD;
mem[16'hBED9] = 8'h85;
mem[16'hBEDA] = 8'h56;
mem[16'hBEDB] = 8'h31;
mem[16'hBEDC] = 8'hCF;
mem[16'hBEDD] = 8'hB8;
mem[16'hBEDE] = 8'h22;
mem[16'hBEDF] = 8'h83;
mem[16'hBEE0] = 8'h5C;
mem[16'hBEE1] = 8'h84;
mem[16'hBEE2] = 8'hC9;
mem[16'hBEE3] = 8'h9F;
mem[16'hBEE4] = 8'h4E;
mem[16'hBEE5] = 8'hEC;
mem[16'hBEE6] = 8'h47;
mem[16'hBEE7] = 8'h02;
mem[16'hBEE8] = 8'h54;
mem[16'hBEE9] = 8'h95;
mem[16'hBEEA] = 8'h40;
mem[16'hBEEB] = 8'hE2;
mem[16'hBEEC] = 8'h4D;
mem[16'hBEED] = 8'h08;
mem[16'hBEEE] = 8'h72;
mem[16'hBEEF] = 8'hC6;
mem[16'hBEF0] = 8'h51;
mem[16'hBEF1] = 8'hF0;
mem[16'hBEF2] = 8'hDF;
mem[16'hBEF3] = 8'h9F;
mem[16'hBEF4] = 8'hF1;
mem[16'hBEF5] = 8'hA1;
mem[16'hBEF6] = 8'h7A;
mem[16'hBEF7] = 8'h1D;
mem[16'hBEF8] = 8'hEB;
mem[16'hBEF9] = 8'h9C;
mem[16'hBEFA] = 8'hC0;
mem[16'hBEFB] = 8'hA7;
mem[16'hBEFC] = 8'h42;
mem[16'hBEFD] = 8'h98;
mem[16'hBEFE] = 8'hEB;
mem[16'hBEFF] = 8'h83;
mem[16'hBF00] = 8'hA4;
mem[16'hBF01] = 8'h08;
mem[16'hBF02] = 8'hA3;
mem[16'hBF03] = 8'hA6;
mem[16'hBF04] = 8'hAC;
mem[16'hBF05] = 8'h2C;
mem[16'hBF06] = 8'hA7;
mem[16'hBF07] = 8'h7B;
mem[16'hBF08] = 8'hA2;
mem[16'hBF09] = 8'h00;
mem[16'hBF0A] = 8'hAB;
mem[16'hBF0B] = 8'hAE;
mem[16'hBF0C] = 8'hAC;
mem[16'hBF0D] = 8'h24;
mem[16'hBF0E] = 8'hAF;
mem[16'hBF0F] = 8'h0A;
mem[16'hBF10] = 8'h4C;
mem[16'hBF11] = 8'h9D;
mem[16'hBF12] = 8'hF8;
mem[16'hBF13] = 8'h00;
mem[16'hBF14] = 8'h71;
mem[16'hBF15] = 8'hE9;
mem[16'hBF16] = 8'h4A;
mem[16'hBF17] = 8'hA9;
mem[16'hBF18] = 8'h7D;
mem[16'hBF19] = 8'h32;
mem[16'hBF1A] = 8'h66;
mem[16'hBF1B] = 8'hBF;
mem[16'hBF1C] = 8'h15;
mem[16'hBF1D] = 8'hBC;
mem[16'hBF1E] = 8'hBB;
mem[16'hBF1F] = 8'hF3;
mem[16'hBF20] = 8'h09;
mem[16'hBF21] = 8'h80;
mem[16'hBF22] = 8'h5E;
mem[16'hBF23] = 8'h89;
mem[16'hBF24] = 8'h2D;
mem[16'hBF25] = 8'h84;
mem[16'hBF26] = 8'h83;
mem[16'hBF27] = 8'h4B;
mem[16'hBF28] = 8'h01;
mem[16'hBF29] = 8'h88;
mem[16'hBF2A] = 8'h23;
mem[16'hBF2B] = 8'h8A;
mem[16'hBF2C] = 8'h0D;
mem[16'hBF2D] = 8'h91;
mem[16'hBF2E] = 8'h22;
mem[16'hBF2F] = 8'h4E;
mem[16'hBF30] = 8'h7C;
mem[16'hBF31] = 8'h29;
mem[16'hBF32] = 8'h6E;
mem[16'hBF33] = 8'h9C;
mem[16'hBF34] = 8'h76;
mem[16'hBF35] = 8'h91;
mem[16'hBF36] = 8'h3A;
mem[16'hBF37] = 8'h36;
mem[16'hBF38] = 8'h9C;
mem[16'hBF39] = 8'h35;
mem[16'hBF3A] = 8'h66;
mem[16'hBF3B] = 8'h93;
mem[16'hBF3C] = 8'hDC;
mem[16'hBF3D] = 8'hE1;
mem[16'hBF3E] = 8'h2D;
mem[16'hBF3F] = 8'h3A;
mem[16'hBF40] = 8'h45;
mem[16'hBF41] = 8'h1D;
mem[16'hBF42] = 8'h63;
mem[16'hBF43] = 8'hD5;
mem[16'hBF44] = 8'h57;
mem[16'hBF45] = 8'h89;
mem[16'hBF46] = 8'h6F;
mem[16'hBF47] = 8'hFA;
mem[16'hBF48] = 8'h44;
mem[16'hBF49] = 8'hE5;
mem[16'hBF4A] = 8'h62;
mem[16'hBF4B] = 8'hF7;
mem[16'hBF4C] = 8'hF8;
mem[16'hBF4D] = 8'h88;
mem[16'hBF4E] = 8'hEA;
mem[16'hBF4F] = 8'h49;
mem[16'hBF50] = 8'h64;
mem[16'hBF51] = 8'hAC;
mem[16'hBF52] = 8'hEE;
mem[16'hBF53] = 8'h37;
mem[16'hBF54] = 8'h28;
mem[16'hBF55] = 8'h02;
mem[16'hBF56] = 8'h1C;
mem[16'hBF57] = 8'hEA;
mem[16'hBF58] = 8'h10;
mem[16'hBF59] = 8'hE4;
mem[16'hBF5A] = 8'h26;
mem[16'hBF5B] = 8'h02;
mem[16'hBF5C] = 8'h90;
mem[16'hBF5D] = 8'hD1;
mem[16'hBF5E] = 8'hF1;
mem[16'hBF5F] = 8'h46;
mem[16'hBF60] = 8'h69;
mem[16'hBF61] = 8'hCB;
mem[16'hBF62] = 8'h1E;
mem[16'hBF63] = 8'hC3;
mem[16'hBF64] = 8'h6C;
mem[16'hBF65] = 8'hD0;
mem[16'hBF66] = 8'h6F;
mem[16'hBF67] = 8'hCB;
mem[16'hBF68] = 8'h49;
mem[16'hBF69] = 8'hC5;
mem[16'hBF6A] = 8'h66;
mem[16'hBF6B] = 8'h5E;
mem[16'hBF6C] = 8'h30;
mem[16'hBF6D] = 8'h75;
mem[16'hBF6E] = 8'hA2;
mem[16'hBF6F] = 8'hDA;
mem[16'hBF70] = 8'h7E;
mem[16'hBF71] = 8'hDC;
mem[16'hBF72] = 8'h44;
mem[16'hBF73] = 8'h51;
mem[16'hBF74] = 8'h2B;
mem[16'hBF75] = 8'hDA;
mem[16'hBF76] = 8'h73;
mem[16'hBF77] = 8'h7B;
mem[16'hBF78] = 8'h74;
mem[16'hBF79] = 8'hD5;
mem[16'hBF7A] = 8'h4F;
mem[16'hBF7B] = 8'hD7;
mem[16'hBF7C] = 8'hD8;
mem[16'hBF7D] = 8'h48;
mem[16'hBF7E] = 8'hD2;
mem[16'hBF7F] = 8'hDA;
mem[16'hBF80] = 8'hB5;
mem[16'hBF81] = 8'h2D;
mem[16'hBF82] = 8'h24;
mem[16'hBF83] = 8'hB6;
mem[16'hBF84] = 8'h28;
mem[16'hBF85] = 8'h22;
mem[16'hBF86] = 8'hE2;
mem[16'hBF87] = 8'hFB;
mem[16'hBF88] = 8'hD5;
mem[16'hBF89] = 8'h85;
mem[16'hBF8A] = 8'h2E;
mem[16'hBF8B] = 8'h9E;
mem[16'hBF8C] = 8'hA6;
mem[16'hBF8D] = 8'h9A;
mem[16'hBF8E] = 8'hBB;
mem[16'hBF8F] = 8'h23;
mem[16'hBF90] = 8'h34;
mem[16'hBF91] = 8'hB5;
mem[16'hBF92] = 8'h2E;
mem[16'hBF93] = 8'hC8;
mem[16'hBF94] = 8'h08;
mem[16'hBF95] = 8'h38;
mem[16'hBF96] = 8'hBF;
mem[16'hBF97] = 8'h9B;
mem[16'hBF98] = 8'h0C;
mem[16'hBF99] = 8'h98;
mem[16'hBF9A] = 8'h63;
mem[16'hBF9B] = 8'hF7;
mem[16'hBF9C] = 8'h9D;
mem[16'hBF9D] = 8'h60;
mem[16'hBF9E] = 8'hF2;
mem[16'hBF9F] = 8'h8A;
mem[16'hBFA0] = 8'hBA;
mem[16'hBFA1] = 8'hB2;
mem[16'hBFA2] = 8'h97;
mem[16'hBFA3] = 8'h0F;
mem[16'hBFA4] = 8'h0C;
mem[16'hBFA5] = 8'h81;
mem[16'hBFA6] = 8'h1A;
mem[16'hBFA7] = 8'hFC;
mem[16'hBFA8] = 8'hA4;
mem[16'hBFA9] = 8'h0A;
mem[16'hBFAA] = 8'hBF;
mem[16'hBFAB] = 8'hE8;
mem[16'hBFAC] = 8'hBF;
mem[16'hBFAD] = 8'h98;
mem[16'hBFAE] = 8'hF2;
mem[16'hBFAF] = 8'h02;
mem[16'hBFB0] = 8'h94;
mem[16'hBFB1] = 8'h0D;
mem[16'hBFB2] = 8'hE9;
mem[16'hBFB3] = 8'h53;
mem[16'hBFB4] = 8'h18;
mem[16'hBFB5] = 8'h1D;
mem[16'hBFB6] = 8'hBA;
mem[16'hBFB7] = 8'h1B;
mem[16'hBFB8] = 8'h90;
mem[16'hBFB9] = 8'h15;
mem[16'hBFBA] = 8'h92;
mem[16'hBFBB] = 8'h16;
mem[16'hBFBC] = 8'hB9;
mem[16'hBFBD] = 8'h11;
mem[16'hBFBE] = 8'hB4;
mem[16'hBFBF] = 8'h12;
mem[16'hBFC0] = 8'h9C;
mem[16'hBFC1] = 8'h6B;
mem[16'hBFC2] = 8'h8E;
mem[16'hBFC3] = 8'h63;
mem[16'hBFC4] = 8'hD8;
mem[16'hBFC5] = 8'h6B;
mem[16'hBFC6] = 8'hC3;
mem[16'hBFC7] = 8'hCB;
mem[16'hBFC8] = 8'hF5;
mem[16'hBFC9] = 8'h65;
mem[16'hBFCA] = 8'hAE;
mem[16'hBFCB] = 8'hB7;
mem[16'hBFCC] = 8'h9B;
mem[16'hBFCD] = 8'h87;
mem[16'hBFCE] = 8'h63;
mem[16'hBFCF] = 8'h93;
mem[16'hBFD0] = 8'h69;
mem[16'hBFD1] = 8'hD8;
mem[16'hBFD2] = 8'h7F;
mem[16'hBFD3] = 8'hB6;
mem[16'hBFD4] = 8'h79;
mem[16'hBFD5] = 8'h89;
mem[16'hBFD6] = 8'h8C;
mem[16'hBFD7] = 8'hB2;
mem[16'hBFD8] = 8'h70;
mem[16'hBFD9] = 8'h85;
mem[16'hBFDA] = 8'h84;
mem[16'hBFDB] = 8'hBE;
mem[16'hBFDC] = 8'h78;
mem[16'hBFDD] = 8'h81;
mem[16'hBFDE] = 8'h9C;
mem[16'hBFDF] = 8'hBA;
mem[16'hBFE0] = 8'h8C;
mem[16'hBFE1] = 8'hBD;
mem[16'hBFE2] = 8'hA4;
mem[16'hBFE3] = 8'h9F;
mem[16'hBFE4] = 8'h9F;
mem[16'hBFE5] = 8'hE0;
mem[16'hBFE6] = 8'hE7;
mem[16'hBFE7] = 8'hCA;
mem[16'hBFE8] = 8'h84;
mem[16'hBFE9] = 8'hE8;
mem[16'hBFEA] = 8'h17;
mem[16'hBFEB] = 8'h87;
mem[16'hBFEC] = 8'h0C;
mem[16'hBFED] = 8'hB1;
mem[16'hBFEE] = 8'h43;
mem[16'hBFEF] = 8'hE3;
mem[16'hBFF0] = 8'h5C;
mem[16'hBFF1] = 8'hF4;
mem[16'hBFF2] = 8'hFE;
mem[16'hBFF3] = 8'hC6;
mem[16'hBFF4] = 8'h58;
mem[16'hBFF5] = 8'h5D;
mem[16'hBFF6] = 8'h92;
mem[16'hBFF7] = 8'h8B;
mem[16'hBFF8] = 8'hAE;
mem[16'hBFF9] = 8'hF8;
mem[16'hBFFA] = 8'h02;
mem[16'hBFFB] = 8'h97;
mem[16'hBFFC] = 8'h3C;
mem[16'hBFFD] = 8'hAD;
mem[16'hBFFE] = 8'hAD;
mem[16'hBFFF] = 8'h53;
mem[16'hC000] = 8'h00;
mem[16'hC001] = 8'h00;
mem[16'hC002] = 8'h00;
mem[16'hC003] = 8'h00;
mem[16'hC004] = 8'h00;
mem[16'hC005] = 8'h00;
mem[16'hC006] = 8'h00;
mem[16'hC007] = 8'h00;
mem[16'hC008] = 8'h00;
mem[16'hC009] = 8'h00;
mem[16'hC00A] = 8'h00;
mem[16'hC00B] = 8'h00;
mem[16'hC00C] = 8'h00;
mem[16'hC00D] = 8'h00;
mem[16'hC00E] = 8'h00;
mem[16'hC00F] = 8'h00;
mem[16'hC010] = 8'h00;
mem[16'hC011] = 8'h00;
mem[16'hC012] = 8'h00;
mem[16'hC013] = 8'h00;
mem[16'hC014] = 8'h00;
mem[16'hC015] = 8'h00;
mem[16'hC016] = 8'h00;
mem[16'hC017] = 8'h00;
mem[16'hC018] = 8'h00;
mem[16'hC019] = 8'h00;
mem[16'hC01A] = 8'h00;
mem[16'hC01B] = 8'h00;
mem[16'hC01C] = 8'h00;
mem[16'hC01D] = 8'h00;
mem[16'hC01E] = 8'h00;
mem[16'hC01F] = 8'h00;
mem[16'hC020] = 8'h00;
mem[16'hC021] = 8'h00;
mem[16'hC022] = 8'h00;
mem[16'hC023] = 8'h00;
mem[16'hC024] = 8'h00;
mem[16'hC025] = 8'h00;
mem[16'hC026] = 8'h00;
mem[16'hC027] = 8'h00;
mem[16'hC028] = 8'h00;
mem[16'hC029] = 8'h00;
mem[16'hC02A] = 8'h00;
mem[16'hC02B] = 8'h00;
mem[16'hC02C] = 8'h00;
mem[16'hC02D] = 8'h00;
mem[16'hC02E] = 8'h00;
mem[16'hC02F] = 8'h00;
mem[16'hC030] = 8'h00;
mem[16'hC031] = 8'h00;
mem[16'hC032] = 8'h00;
mem[16'hC033] = 8'h00;
mem[16'hC034] = 8'h00;
mem[16'hC035] = 8'h00;
mem[16'hC036] = 8'h00;
mem[16'hC037] = 8'h00;
mem[16'hC038] = 8'h00;
mem[16'hC039] = 8'h00;
mem[16'hC03A] = 8'h00;
mem[16'hC03B] = 8'h00;
mem[16'hC03C] = 8'h00;
mem[16'hC03D] = 8'h00;
mem[16'hC03E] = 8'h00;
mem[16'hC03F] = 8'h00;
mem[16'hC040] = 8'h00;
mem[16'hC041] = 8'h00;
mem[16'hC042] = 8'h00;
mem[16'hC043] = 8'h00;
mem[16'hC044] = 8'h00;
mem[16'hC045] = 8'h00;
mem[16'hC046] = 8'h00;
mem[16'hC047] = 8'h00;
mem[16'hC048] = 8'h00;
mem[16'hC049] = 8'h00;
mem[16'hC04A] = 8'h00;
mem[16'hC04B] = 8'h00;
mem[16'hC04C] = 8'h00;
mem[16'hC04D] = 8'h00;
mem[16'hC04E] = 8'h00;
mem[16'hC04F] = 8'h00;
mem[16'hC050] = 8'h00;
mem[16'hC051] = 8'h00;
mem[16'hC052] = 8'h00;
mem[16'hC053] = 8'h00;
mem[16'hC054] = 8'h00;
mem[16'hC055] = 8'h00;
mem[16'hC056] = 8'h00;
mem[16'hC057] = 8'h00;
mem[16'hC058] = 8'h00;
mem[16'hC059] = 8'h00;
mem[16'hC05A] = 8'h00;
mem[16'hC05B] = 8'h00;
mem[16'hC05C] = 8'h00;
mem[16'hC05D] = 8'h00;
mem[16'hC05E] = 8'h00;
mem[16'hC05F] = 8'h00;
mem[16'hC060] = 8'h00;
mem[16'hC061] = 8'h00;
mem[16'hC062] = 8'h00;
mem[16'hC063] = 8'h00;
mem[16'hC064] = 8'h00;
mem[16'hC065] = 8'h00;
mem[16'hC066] = 8'h00;
mem[16'hC067] = 8'h00;
mem[16'hC068] = 8'h00;
mem[16'hC069] = 8'h00;
mem[16'hC06A] = 8'h00;
mem[16'hC06B] = 8'h00;
mem[16'hC06C] = 8'h00;
mem[16'hC06D] = 8'h00;
mem[16'hC06E] = 8'h00;
mem[16'hC06F] = 8'h00;
mem[16'hC070] = 8'h00;
mem[16'hC071] = 8'h00;
mem[16'hC072] = 8'h00;
mem[16'hC073] = 8'h00;
mem[16'hC074] = 8'h00;
mem[16'hC075] = 8'h00;
mem[16'hC076] = 8'h00;
mem[16'hC077] = 8'h00;
mem[16'hC078] = 8'h00;
mem[16'hC079] = 8'h00;
mem[16'hC07A] = 8'h00;
mem[16'hC07B] = 8'h00;
mem[16'hC07C] = 8'h00;
mem[16'hC07D] = 8'h00;
mem[16'hC07E] = 8'h00;
mem[16'hC07F] = 8'h00;
mem[16'hC080] = 8'h00;
mem[16'hC081] = 8'h00;
mem[16'hC082] = 8'h00;
mem[16'hC083] = 8'h00;
mem[16'hC084] = 8'h00;
mem[16'hC085] = 8'h00;
mem[16'hC086] = 8'h00;
mem[16'hC087] = 8'h00;
mem[16'hC088] = 8'h00;
mem[16'hC089] = 8'h00;
mem[16'hC08A] = 8'h00;
mem[16'hC08B] = 8'h00;
mem[16'hC08C] = 8'h00;
mem[16'hC08D] = 8'h00;
mem[16'hC08E] = 8'h00;
mem[16'hC08F] = 8'h00;
mem[16'hC090] = 8'h00;
mem[16'hC091] = 8'h00;
mem[16'hC092] = 8'h00;
mem[16'hC093] = 8'h00;
mem[16'hC094] = 8'h00;
mem[16'hC095] = 8'h00;
mem[16'hC096] = 8'h00;
mem[16'hC097] = 8'h00;
mem[16'hC098] = 8'h00;
mem[16'hC099] = 8'h00;
mem[16'hC09A] = 8'h00;
mem[16'hC09B] = 8'h00;
mem[16'hC09C] = 8'h00;
mem[16'hC09D] = 8'h00;
mem[16'hC09E] = 8'h00;
mem[16'hC09F] = 8'h00;
mem[16'hC0A0] = 8'h00;
mem[16'hC0A1] = 8'h00;
mem[16'hC0A2] = 8'h00;
mem[16'hC0A3] = 8'h00;
mem[16'hC0A4] = 8'h00;
mem[16'hC0A5] = 8'h00;
mem[16'hC0A6] = 8'h00;
mem[16'hC0A7] = 8'h00;
mem[16'hC0A8] = 8'h00;
mem[16'hC0A9] = 8'h00;
mem[16'hC0AA] = 8'h00;
mem[16'hC0AB] = 8'h00;
mem[16'hC0AC] = 8'h00;
mem[16'hC0AD] = 8'h00;
mem[16'hC0AE] = 8'h00;
mem[16'hC0AF] = 8'h00;
mem[16'hC0B0] = 8'h00;
mem[16'hC0B1] = 8'h00;
mem[16'hC0B2] = 8'h00;
mem[16'hC0B3] = 8'h00;
mem[16'hC0B4] = 8'h00;
mem[16'hC0B5] = 8'h00;
mem[16'hC0B6] = 8'h00;
mem[16'hC0B7] = 8'h00;
mem[16'hC0B8] = 8'h00;
mem[16'hC0B9] = 8'h00;
mem[16'hC0BA] = 8'h00;
mem[16'hC0BB] = 8'h00;
mem[16'hC0BC] = 8'h00;
mem[16'hC0BD] = 8'h00;
mem[16'hC0BE] = 8'h00;
mem[16'hC0BF] = 8'h00;
mem[16'hC0C0] = 8'h00;
mem[16'hC0C1] = 8'h00;
mem[16'hC0C2] = 8'h00;
mem[16'hC0C3] = 8'h00;
mem[16'hC0C4] = 8'h00;
mem[16'hC0C5] = 8'h00;
mem[16'hC0C6] = 8'h00;
mem[16'hC0C7] = 8'h00;
mem[16'hC0C8] = 8'h00;
mem[16'hC0C9] = 8'h00;
mem[16'hC0CA] = 8'h00;
mem[16'hC0CB] = 8'h00;
mem[16'hC0CC] = 8'h00;
mem[16'hC0CD] = 8'h00;
mem[16'hC0CE] = 8'h00;
mem[16'hC0CF] = 8'h00;
mem[16'hC0D0] = 8'h00;
mem[16'hC0D1] = 8'h00;
mem[16'hC0D2] = 8'h00;
mem[16'hC0D3] = 8'h00;
mem[16'hC0D4] = 8'h00;
mem[16'hC0D5] = 8'h00;
mem[16'hC0D6] = 8'h00;
mem[16'hC0D7] = 8'h00;
mem[16'hC0D8] = 8'h00;
mem[16'hC0D9] = 8'h00;
mem[16'hC0DA] = 8'h00;
mem[16'hC0DB] = 8'h00;
mem[16'hC0DC] = 8'h00;
mem[16'hC0DD] = 8'h00;
mem[16'hC0DE] = 8'h00;
mem[16'hC0DF] = 8'h00;
mem[16'hC0E0] = 8'h00;
mem[16'hC0E1] = 8'h00;
mem[16'hC0E2] = 8'h00;
mem[16'hC0E3] = 8'h00;
mem[16'hC0E4] = 8'h00;
mem[16'hC0E5] = 8'h00;
mem[16'hC0E6] = 8'h00;
mem[16'hC0E7] = 8'h00;
mem[16'hC0E8] = 8'h00;
mem[16'hC0E9] = 8'h00;
mem[16'hC0EA] = 8'h00;
mem[16'hC0EB] = 8'h00;
mem[16'hC0EC] = 8'h00;
mem[16'hC0ED] = 8'h00;
mem[16'hC0EE] = 8'h00;
mem[16'hC0EF] = 8'h00;
mem[16'hC0F0] = 8'h00;
mem[16'hC0F1] = 8'h00;
mem[16'hC0F2] = 8'h00;
mem[16'hC0F3] = 8'h00;
mem[16'hC0F4] = 8'h00;
mem[16'hC0F5] = 8'h00;
mem[16'hC0F6] = 8'h00;
mem[16'hC0F7] = 8'h00;
mem[16'hC0F8] = 8'h00;
mem[16'hC0F9] = 8'h00;
mem[16'hC0FA] = 8'h00;
mem[16'hC0FB] = 8'h00;
mem[16'hC0FC] = 8'h00;
mem[16'hC0FD] = 8'h00;
mem[16'hC0FE] = 8'h00;
mem[16'hC0FF] = 8'h00;
mem[16'hC100] = 8'h18;
mem[16'hC101] = 8'hB0;
mem[16'hC102] = 8'h38;
mem[16'hC103] = 8'h48;
mem[16'hC104] = 8'h8A;
mem[16'hC105] = 8'h48;
mem[16'hC106] = 8'h98;
mem[16'hC107] = 8'h48;
mem[16'hC108] = 8'h08;
mem[16'hC109] = 8'h78;
mem[16'hC10A] = 8'h20;
mem[16'hC10B] = 8'h58;
mem[16'hC10C] = 8'hFF;
mem[16'hC10D] = 8'hBA;
mem[16'hC10E] = 8'h68;
mem[16'hC10F] = 8'h68;
mem[16'hC110] = 8'h68;
mem[16'hC111] = 8'h68;
mem[16'hC112] = 8'hA8;
mem[16'hC113] = 8'hCA;
mem[16'hC114] = 8'h9A;
mem[16'hC115] = 8'h68;
mem[16'hC116] = 8'h28;
mem[16'hC117] = 8'hAA;
mem[16'hC118] = 8'h90;
mem[16'hC119] = 8'h38;
mem[16'hC11A] = 8'hBD;
mem[16'hC11B] = 8'hB8;
mem[16'hC11C] = 8'h05;
mem[16'hC11D] = 8'h10;
mem[16'hC11E] = 8'h19;
mem[16'hC11F] = 8'h98;
mem[16'hC120] = 8'h29;
mem[16'hC121] = 8'h7F;
mem[16'hC122] = 8'h49;
mem[16'hC123] = 8'h30;
mem[16'hC124] = 8'hC9;
mem[16'hC125] = 8'h0A;
mem[16'hC126] = 8'h90;
mem[16'hC127] = 8'h3B;
mem[16'hC128] = 8'hC9;
mem[16'hC129] = 8'h78;
mem[16'hC12A] = 8'hB0;
mem[16'hC12B] = 8'h29;
mem[16'hC12C] = 8'h49;
mem[16'hC12D] = 8'h3D;
mem[16'hC12E] = 8'hF0;
mem[16'hC12F] = 8'h21;
mem[16'hC130] = 8'h98;
mem[16'hC131] = 8'h29;
mem[16'hC132] = 8'h9F;
mem[16'hC133] = 8'h9D;
mem[16'hC134] = 8'h38;
mem[16'hC135] = 8'h06;
mem[16'hC136] = 8'h90;
mem[16'hC137] = 8'h7E;
mem[16'hC138] = 8'hBD;
mem[16'hC139] = 8'hB8;
mem[16'hC13A] = 8'h06;
mem[16'hC13B] = 8'h30;
mem[16'hC13C] = 8'h14;
mem[16'hC13D] = 8'hA5;
mem[16'hC13E] = 8'h24;
mem[16'hC13F] = 8'hDD;
mem[16'hC140] = 8'h38;
mem[16'hC141] = 8'h07;
mem[16'hC142] = 8'hB0;
mem[16'hC143] = 8'h0D;
mem[16'hC144] = 8'hC9;
mem[16'hC145] = 8'h11;
mem[16'hC146] = 8'hB0;
mem[16'hC147] = 8'h09;
mem[16'hC148] = 8'h09;
mem[16'hC149] = 8'hF0;
mem[16'hC14A] = 8'h3D;
mem[16'hC14B] = 8'h38;
mem[16'hC14C] = 8'h07;
mem[16'hC14D] = 8'h65;
mem[16'hC14E] = 8'h24;
mem[16'hC14F] = 8'h85;
mem[16'hC150] = 8'h24;
mem[16'hC151] = 8'h4A;
mem[16'hC152] = 8'h38;
mem[16'hC153] = 8'hB0;
mem[16'hC154] = 8'h6D;
mem[16'hC155] = 8'h18;
mem[16'hC156] = 8'h6A;
mem[16'hC157] = 8'h3D;
mem[16'hC158] = 8'hB8;
mem[16'hC159] = 8'h06;
mem[16'hC15A] = 8'h90;
mem[16'hC15B] = 8'h02;
mem[16'hC15C] = 8'h49;
mem[16'hC15D] = 8'h81;
mem[16'hC15E] = 8'h9D;
mem[16'hC15F] = 8'hB8;
mem[16'hC160] = 8'h06;
mem[16'hC161] = 8'hD0;
mem[16'hC162] = 8'h53;
mem[16'hC163] = 8'hA0;
mem[16'hC164] = 8'h0A;
mem[16'hC165] = 8'h7D;
mem[16'hC166] = 8'h38;
mem[16'hC167] = 8'h05;
mem[16'hC168] = 8'h88;
mem[16'hC169] = 8'hD0;
mem[16'hC16A] = 8'hFA;
mem[16'hC16B] = 8'h9D;
mem[16'hC16C] = 8'hB8;
mem[16'hC16D] = 8'h04;
mem[16'hC16E] = 8'h9D;
mem[16'hC16F] = 8'h38;
mem[16'hC170] = 8'h05;
mem[16'hC171] = 8'h38;
mem[16'hC172] = 8'hB0;
mem[16'hC173] = 8'h43;
mem[16'hC174] = 8'hC5;
mem[16'hC175] = 8'h24;
mem[16'hC176] = 8'h90;
mem[16'hC177] = 8'h3A;
mem[16'hC178] = 8'h68;
mem[16'hC179] = 8'hA8;
mem[16'hC17A] = 8'h68;
mem[16'hC17B] = 8'hAA;
mem[16'hC17C] = 8'h68;
mem[16'hC17D] = 8'h4C;
mem[16'hC17E] = 8'hF0;
mem[16'hC17F] = 8'hFD;
mem[16'hC180] = 8'h90;
mem[16'hC181] = 8'hFE;
mem[16'hC182] = 8'hB0;
mem[16'hC183] = 8'hFE;
mem[16'hC184] = 8'h99;
mem[16'hC185] = 8'h80;
mem[16'hC186] = 8'hC0;
mem[16'hC187] = 8'h90;
mem[16'hC188] = 8'h37;
mem[16'hC189] = 8'h49;
mem[16'hC18A] = 8'h07;
mem[16'hC18B] = 8'hA8;
mem[16'hC18C] = 8'h49;
mem[16'hC18D] = 8'h0A;
mem[16'hC18E] = 8'h0A;
mem[16'hC18F] = 8'hD0;
mem[16'hC190] = 8'h06;
mem[16'hC191] = 8'hB8;
mem[16'hC192] = 8'h85;
mem[16'hC193] = 8'h24;
mem[16'hC194] = 8'h9D;
mem[16'hC195] = 8'h38;
mem[16'hC196] = 8'h07;
mem[16'hC197] = 8'hBD;
mem[16'hC198] = 8'hB8;
mem[16'hC199] = 8'h06;
mem[16'hC19A] = 8'h4A;
mem[16'hC19B] = 8'h70;
mem[16'hC19C] = 8'h02;
mem[16'hC19D] = 8'hB0;
mem[16'hC19E] = 8'h23;
mem[16'hC19F] = 8'h0A;
mem[16'hC1A0] = 8'h0A;
mem[16'hC1A1] = 8'hA9;
mem[16'hC1A2] = 8'h27;
mem[16'hC1A3] = 8'hB0;
mem[16'hC1A4] = 8'hCF;
mem[16'hC1A5] = 8'hBD;
mem[16'hC1A6] = 8'h38;
mem[16'hC1A7] = 8'h07;
mem[16'hC1A8] = 8'hFD;
mem[16'hC1A9] = 8'hB8;
mem[16'hC1AA] = 8'h04;
mem[16'hC1AB] = 8'hC9;
mem[16'hC1AC] = 8'hF8;
mem[16'hC1AD] = 8'h90;
mem[16'hC1AE] = 8'h03;
mem[16'hC1AF] = 8'h69;
mem[16'hC1B0] = 8'h27;
mem[16'hC1B1] = 8'hAC;
mem[16'hC1B2] = 8'hA9;
mem[16'hC1B3] = 8'h00;
mem[16'hC1B4] = 8'h85;
mem[16'hC1B5] = 8'h24;
mem[16'hC1B6] = 8'h18;
mem[16'hC1B7] = 8'h7E;
mem[16'hC1B8] = 8'hB8;
mem[16'hC1B9] = 8'h05;
mem[16'hC1BA] = 8'h68;
mem[16'hC1BB] = 8'hA8;
mem[16'hC1BC] = 8'h68;
mem[16'hC1BD] = 8'hAA;
mem[16'hC1BE] = 8'h68;
mem[16'hC1BF] = 8'h60;
mem[16'hC1C0] = 8'h90;
mem[16'hC1C1] = 8'h27;
mem[16'hC1C2] = 8'hB0;
mem[16'hC1C3] = 8'h00;
mem[16'hC1C4] = 8'h10;
mem[16'hC1C5] = 8'h11;
mem[16'hC1C6] = 8'hA9;
mem[16'hC1C7] = 8'h89;
mem[16'hC1C8] = 8'h9D;
mem[16'hC1C9] = 8'h38;
mem[16'hC1CA] = 8'h06;
mem[16'hC1CB] = 8'h9D;
mem[16'hC1CC] = 8'hB8;
mem[16'hC1CD] = 8'h06;
mem[16'hC1CE] = 8'hA9;
mem[16'hC1CF] = 8'h28;
mem[16'hC1D0] = 8'h9D;
mem[16'hC1D1] = 8'hB8;
mem[16'hC1D2] = 8'h04;
mem[16'hC1D3] = 8'hA9;
mem[16'hC1D4] = 8'h02;
mem[16'hC1D5] = 8'h85;
mem[16'hC1D6] = 8'h36;
mem[16'hC1D7] = 8'h98;
mem[16'hC1D8] = 8'h5D;
mem[16'hC1D9] = 8'h38;
mem[16'hC1DA] = 8'h06;
mem[16'hC1DB] = 8'h0A;
mem[16'hC1DC] = 8'hF0;
mem[16'hC1DD] = 8'h90;
mem[16'hC1DE] = 8'h5E;
mem[16'hC1DF] = 8'hB8;
mem[16'hC1E0] = 8'h05;
mem[16'hC1E1] = 8'h98;
mem[16'hC1E2] = 8'h48;
mem[16'hC1E3] = 8'h8A;
mem[16'hC1E4] = 8'h0A;
mem[16'hC1E5] = 8'h0A;
mem[16'hC1E6] = 8'h0A;
mem[16'hC1E7] = 8'h0A;
mem[16'hC1E8] = 8'hA8;
mem[16'hC1E9] = 8'hBD;
mem[16'hC1EA] = 8'h38;
mem[16'hC1EB] = 8'h07;
mem[16'hC1EC] = 8'hC5;
mem[16'hC1ED] = 8'h24;
mem[16'hC1EE] = 8'h68;
mem[16'hC1EF] = 8'hB0;
mem[16'hC1F0] = 8'h05;
mem[16'hC1F1] = 8'h48;
mem[16'hC1F2] = 8'h29;
mem[16'hC1F3] = 8'h80;
mem[16'hC1F4] = 8'h09;
mem[16'hC1F5] = 8'h20;
mem[16'hC1F6] = 8'h2C;
mem[16'hC1F7] = 8'h58;
mem[16'hC1F8] = 8'hFF;
mem[16'hC1F9] = 8'hF0;
mem[16'hC1FA] = 8'h03;
mem[16'hC1FB] = 8'hFE;
mem[16'hC1FC] = 8'h38;
mem[16'hC1FD] = 8'h07;
mem[16'hC1FE] = 8'h70;
mem[16'hC1FF] = 8'h84;
mem[16'hC200] = 8'h2C;
mem[16'hC201] = 8'h58;
mem[16'hC202] = 8'hFF;
mem[16'hC203] = 8'h70;
mem[16'hC204] = 8'h0C;
mem[16'hC205] = 8'h38;
mem[16'hC206] = 8'h90;
mem[16'hC207] = 8'h18;
mem[16'hC208] = 8'hB8;
mem[16'hC209] = 8'h50;
mem[16'hC20A] = 8'h06;
mem[16'hC20B] = 8'h01;
mem[16'hC20C] = 8'h31;
mem[16'hC20D] = 8'h8E;
mem[16'hC20E] = 8'h94;
mem[16'hC20F] = 8'h97;
mem[16'hC210] = 8'h9A;
mem[16'hC211] = 8'h85;
mem[16'hC212] = 8'h27;
mem[16'hC213] = 8'h86;
mem[16'hC214] = 8'h35;
mem[16'hC215] = 8'h8A;
mem[16'hC216] = 8'h48;
mem[16'hC217] = 8'h98;
mem[16'hC218] = 8'h48;
mem[16'hC219] = 8'h08;
mem[16'hC21A] = 8'h78;
mem[16'hC21B] = 8'h8D;
mem[16'hC21C] = 8'hFF;
mem[16'hC21D] = 8'hCF;
mem[16'hC21E] = 8'h20;
mem[16'hC21F] = 8'h58;
mem[16'hC220] = 8'hFF;
mem[16'hC221] = 8'hBA;
mem[16'hC222] = 8'hBD;
mem[16'hC223] = 8'h00;
mem[16'hC224] = 8'h01;
mem[16'hC225] = 8'h8D;
mem[16'hC226] = 8'hF8;
mem[16'hC227] = 8'h07;
mem[16'hC228] = 8'hAA;
mem[16'hC229] = 8'h0A;
mem[16'hC22A] = 8'h0A;
mem[16'hC22B] = 8'h0A;
mem[16'hC22C] = 8'h0A;
mem[16'hC22D] = 8'h85;
mem[16'hC22E] = 8'h26;
mem[16'hC22F] = 8'hA8;
mem[16'hC230] = 8'h28;
mem[16'hC231] = 8'h50;
mem[16'hC232] = 8'h29;
mem[16'hC233] = 8'h1E;
mem[16'hC234] = 8'h38;
mem[16'hC235] = 8'h05;
mem[16'hC236] = 8'h5E;
mem[16'hC237] = 8'h38;
mem[16'hC238] = 8'h05;
mem[16'hC239] = 8'hB9;
mem[16'hC23A] = 8'h8A;
mem[16'hC23B] = 8'hC0;
mem[16'hC23C] = 8'h29;
mem[16'hC23D] = 8'h1F;
mem[16'hC23E] = 8'hD0;
mem[16'hC23F] = 8'h05;
mem[16'hC240] = 8'hA9;
mem[16'hC241] = 8'hEF;
mem[16'hC242] = 8'h20;
mem[16'hC243] = 8'h05;
mem[16'hC244] = 8'hC8;
mem[16'hC245] = 8'hE4;
mem[16'hC246] = 8'h37;
mem[16'hC247] = 8'hD0;
mem[16'hC248] = 8'h0B;
mem[16'hC249] = 8'hA9;
mem[16'hC24A] = 8'h07;
mem[16'hC24B] = 8'hC5;
mem[16'hC24C] = 8'h36;
mem[16'hC24D] = 8'hF0;
mem[16'hC24E] = 8'h05;
mem[16'hC24F] = 8'h85;
mem[16'hC250] = 8'h36;
mem[16'hC251] = 8'h18;
mem[16'hC252] = 8'h90;
mem[16'hC253] = 8'h08;
mem[16'hC254] = 8'hE4;
mem[16'hC255] = 8'h39;
mem[16'hC256] = 8'hD0;
mem[16'hC257] = 8'hF9;
mem[16'hC258] = 8'hA9;
mem[16'hC259] = 8'h05;
mem[16'hC25A] = 8'h85;
mem[16'hC25B] = 8'h38;
mem[16'hC25C] = 8'hBD;
mem[16'hC25D] = 8'h38;
mem[16'hC25E] = 8'h07;
mem[16'hC25F] = 8'h29;
mem[16'hC260] = 8'h02;
mem[16'hC261] = 8'h08;
mem[16'hC262] = 8'h90;
mem[16'hC263] = 8'h03;
mem[16'hC264] = 8'h4C;
mem[16'hC265] = 8'hBF;
mem[16'hC266] = 8'hC8;
mem[16'hC267] = 8'hBD;
mem[16'hC268] = 8'hB8;
mem[16'hC269] = 8'h04;
mem[16'hC26A] = 8'h48;
mem[16'hC26B] = 8'h0A;
mem[16'hC26C] = 8'h10;
mem[16'hC26D] = 8'h0E;
mem[16'hC26E] = 8'hA6;
mem[16'hC26F] = 8'h35;
mem[16'hC270] = 8'hA5;
mem[16'hC271] = 8'h27;
mem[16'hC272] = 8'h09;
mem[16'hC273] = 8'h20;
mem[16'hC274] = 8'h9D;
mem[16'hC275] = 8'h00;
mem[16'hC276] = 8'h02;
mem[16'hC277] = 8'h85;
mem[16'hC278] = 8'h27;
mem[16'hC279] = 8'hAE;
mem[16'hC27A] = 8'hF8;
mem[16'hC27B] = 8'h07;
mem[16'hC27C] = 8'h68;
mem[16'hC27D] = 8'h29;
mem[16'hC27E] = 8'hBF;
mem[16'hC27F] = 8'h9D;
mem[16'hC280] = 8'hB8;
mem[16'hC281] = 8'h04;
mem[16'hC282] = 8'h28;
mem[16'hC283] = 8'hF0;
mem[16'hC284] = 8'h06;
mem[16'hC285] = 8'h20;
mem[16'hC286] = 8'h63;
mem[16'hC287] = 8'hCB;
mem[16'hC288] = 8'h4C;
mem[16'hC289] = 8'hB5;
mem[16'hC28A] = 8'hC8;
mem[16'hC28B] = 8'h4C;
mem[16'hC28C] = 8'hFC;
mem[16'hC28D] = 8'hC8;
mem[16'hC28E] = 8'h20;
mem[16'hC28F] = 8'h00;
mem[16'hC290] = 8'hC8;
mem[16'hC291] = 8'hA2;
mem[16'hC292] = 8'h00;
mem[16'hC293] = 8'h60;
mem[16'hC294] = 8'h4C;
mem[16'hC295] = 8'h9B;
mem[16'hC296] = 8'hC8;
mem[16'hC297] = 8'h4C;
mem[16'hC298] = 8'hAA;
mem[16'hC299] = 8'hC9;
mem[16'hC29A] = 8'h4A;
mem[16'hC29B] = 8'h20;
mem[16'hC29C] = 8'h9B;
mem[16'hC29D] = 8'hC9;
mem[16'hC29E] = 8'hB0;
mem[16'hC29F] = 8'h08;
mem[16'hC2A0] = 8'h20;
mem[16'hC2A1] = 8'hF5;
mem[16'hC2A2] = 8'hCA;
mem[16'hC2A3] = 8'hF0;
mem[16'hC2A4] = 8'h06;
mem[16'hC2A5] = 8'h18;
mem[16'hC2A6] = 8'h90;
mem[16'hC2A7] = 8'h03;
mem[16'hC2A8] = 8'h20;
mem[16'hC2A9] = 8'hD2;
mem[16'hC2AA] = 8'hCA;
mem[16'hC2AB] = 8'hBD;
mem[16'hC2AC] = 8'hB8;
mem[16'hC2AD] = 8'h05;
mem[16'hC2AE] = 8'hAA;
mem[16'hC2AF] = 8'h60;
mem[16'hC2B0] = 8'hA2;
mem[16'hC2B1] = 8'h03;
mem[16'hC2B2] = 8'hB5;
mem[16'hC2B3] = 8'h36;
mem[16'hC2B4] = 8'h48;
mem[16'hC2B5] = 8'hCA;
mem[16'hC2B6] = 8'h10;
mem[16'hC2B7] = 8'hFA;
mem[16'hC2B8] = 8'hAE;
mem[16'hC2B9] = 8'hF8;
mem[16'hC2BA] = 8'h07;
mem[16'hC2BB] = 8'hBD;
mem[16'hC2BC] = 8'h38;
mem[16'hC2BD] = 8'h06;
mem[16'hC2BE] = 8'h85;
mem[16'hC2BF] = 8'h36;
mem[16'hC2C0] = 8'hBD;
mem[16'hC2C1] = 8'hB8;
mem[16'hC2C2] = 8'h04;
mem[16'hC2C3] = 8'h29;
mem[16'hC2C4] = 8'h38;
mem[16'hC2C5] = 8'h4A;
mem[16'hC2C6] = 8'h4A;
mem[16'hC2C7] = 8'h4A;
mem[16'hC2C8] = 8'h09;
mem[16'hC2C9] = 8'hC0;
mem[16'hC2CA] = 8'h85;
mem[16'hC2CB] = 8'h37;
mem[16'hC2CC] = 8'h8A;
mem[16'hC2CD] = 8'h48;
mem[16'hC2CE] = 8'hA5;
mem[16'hC2CF] = 8'h27;
mem[16'hC2D0] = 8'h48;
mem[16'hC2D1] = 8'h09;
mem[16'hC2D2] = 8'h80;
mem[16'hC2D3] = 8'h20;
mem[16'hC2D4] = 8'hED;
mem[16'hC2D5] = 8'hFD;
mem[16'hC2D6] = 8'h68;
mem[16'hC2D7] = 8'h85;
mem[16'hC2D8] = 8'h27;
mem[16'hC2D9] = 8'h68;
mem[16'hC2DA] = 8'h8D;
mem[16'hC2DB] = 8'hF8;
mem[16'hC2DC] = 8'h07;
mem[16'hC2DD] = 8'hAA;
mem[16'hC2DE] = 8'h0A;
mem[16'hC2DF] = 8'h0A;
mem[16'hC2E0] = 8'h0A;
mem[16'hC2E1] = 8'h0A;
mem[16'hC2E2] = 8'h85;
mem[16'hC2E3] = 8'h26;
mem[16'hC2E4] = 8'h8D;
mem[16'hC2E5] = 8'hFF;
mem[16'hC2E6] = 8'hCF;
mem[16'hC2E7] = 8'hA5;
mem[16'hC2E8] = 8'h36;
mem[16'hC2E9] = 8'h9D;
mem[16'hC2EA] = 8'h38;
mem[16'hC2EB] = 8'h06;
mem[16'hC2EC] = 8'hA2;
mem[16'hC2ED] = 8'h00;
mem[16'hC2EE] = 8'h68;
mem[16'hC2EF] = 8'h95;
mem[16'hC2F0] = 8'h36;
mem[16'hC2F1] = 8'hE8;
mem[16'hC2F2] = 8'hE0;
mem[16'hC2F3] = 8'h04;
mem[16'hC2F4] = 8'h90;
mem[16'hC2F5] = 8'hF8;
mem[16'hC2F6] = 8'hAE;
mem[16'hC2F7] = 8'hF8;
mem[16'hC2F8] = 8'h07;
mem[16'hC2F9] = 8'h60;
mem[16'hC2FA] = 8'hC1;
mem[16'hC2FB] = 8'hD0;
mem[16'hC2FC] = 8'hD0;
mem[16'hC2FD] = 8'hCC;
mem[16'hC2FE] = 8'hC5;
mem[16'hC2FF] = 8'h08;
mem[16'hC300] = 8'h00;
mem[16'hC301] = 8'h00;
mem[16'hC302] = 8'h00;
mem[16'hC303] = 8'h00;
mem[16'hC304] = 8'h00;
mem[16'hC305] = 8'h00;
mem[16'hC306] = 8'h00;
mem[16'hC307] = 8'h00;
mem[16'hC308] = 8'h00;
mem[16'hC309] = 8'h00;
mem[16'hC30A] = 8'h00;
mem[16'hC30B] = 8'h00;
mem[16'hC30C] = 8'h00;
mem[16'hC30D] = 8'h00;
mem[16'hC30E] = 8'h00;
mem[16'hC30F] = 8'h00;
mem[16'hC310] = 8'h00;
mem[16'hC311] = 8'h00;
mem[16'hC312] = 8'h00;
mem[16'hC313] = 8'h00;
mem[16'hC314] = 8'h00;
mem[16'hC315] = 8'h00;
mem[16'hC316] = 8'h00;
mem[16'hC317] = 8'h00;
mem[16'hC318] = 8'h00;
mem[16'hC319] = 8'h00;
mem[16'hC31A] = 8'h00;
mem[16'hC31B] = 8'h00;
mem[16'hC31C] = 8'h00;
mem[16'hC31D] = 8'h00;
mem[16'hC31E] = 8'h00;
mem[16'hC31F] = 8'h00;
mem[16'hC320] = 8'h00;
mem[16'hC321] = 8'h00;
mem[16'hC322] = 8'h00;
mem[16'hC323] = 8'h00;
mem[16'hC324] = 8'h00;
mem[16'hC325] = 8'h00;
mem[16'hC326] = 8'h00;
mem[16'hC327] = 8'h00;
mem[16'hC328] = 8'h00;
mem[16'hC329] = 8'h00;
mem[16'hC32A] = 8'h00;
mem[16'hC32B] = 8'h00;
mem[16'hC32C] = 8'h00;
mem[16'hC32D] = 8'h00;
mem[16'hC32E] = 8'h00;
mem[16'hC32F] = 8'h00;
mem[16'hC330] = 8'h00;
mem[16'hC331] = 8'h00;
mem[16'hC332] = 8'h00;
mem[16'hC333] = 8'h00;
mem[16'hC334] = 8'h00;
mem[16'hC335] = 8'h00;
mem[16'hC336] = 8'h00;
mem[16'hC337] = 8'h00;
mem[16'hC338] = 8'h00;
mem[16'hC339] = 8'h00;
mem[16'hC33A] = 8'h00;
mem[16'hC33B] = 8'h00;
mem[16'hC33C] = 8'h00;
mem[16'hC33D] = 8'h00;
mem[16'hC33E] = 8'h00;
mem[16'hC33F] = 8'h00;
mem[16'hC340] = 8'h00;
mem[16'hC341] = 8'h00;
mem[16'hC342] = 8'h00;
mem[16'hC343] = 8'h00;
mem[16'hC344] = 8'h00;
mem[16'hC345] = 8'h00;
mem[16'hC346] = 8'h00;
mem[16'hC347] = 8'h00;
mem[16'hC348] = 8'h00;
mem[16'hC349] = 8'h00;
mem[16'hC34A] = 8'h00;
mem[16'hC34B] = 8'h00;
mem[16'hC34C] = 8'h00;
mem[16'hC34D] = 8'h00;
mem[16'hC34E] = 8'h00;
mem[16'hC34F] = 8'h00;
mem[16'hC350] = 8'h00;
mem[16'hC351] = 8'h00;
mem[16'hC352] = 8'h00;
mem[16'hC353] = 8'h00;
mem[16'hC354] = 8'h00;
mem[16'hC355] = 8'h00;
mem[16'hC356] = 8'h00;
mem[16'hC357] = 8'h00;
mem[16'hC358] = 8'h00;
mem[16'hC359] = 8'h00;
mem[16'hC35A] = 8'h00;
mem[16'hC35B] = 8'h00;
mem[16'hC35C] = 8'h00;
mem[16'hC35D] = 8'h00;
mem[16'hC35E] = 8'h00;
mem[16'hC35F] = 8'h00;
mem[16'hC360] = 8'h00;
mem[16'hC361] = 8'h00;
mem[16'hC362] = 8'h00;
mem[16'hC363] = 8'h00;
mem[16'hC364] = 8'h00;
mem[16'hC365] = 8'h00;
mem[16'hC366] = 8'h00;
mem[16'hC367] = 8'h00;
mem[16'hC368] = 8'h00;
mem[16'hC369] = 8'h00;
mem[16'hC36A] = 8'h00;
mem[16'hC36B] = 8'h00;
mem[16'hC36C] = 8'h00;
mem[16'hC36D] = 8'h00;
mem[16'hC36E] = 8'h00;
mem[16'hC36F] = 8'h00;
mem[16'hC370] = 8'h00;
mem[16'hC371] = 8'h00;
mem[16'hC372] = 8'h00;
mem[16'hC373] = 8'h00;
mem[16'hC374] = 8'h00;
mem[16'hC375] = 8'h00;
mem[16'hC376] = 8'h00;
mem[16'hC377] = 8'h00;
mem[16'hC378] = 8'h00;
mem[16'hC379] = 8'h00;
mem[16'hC37A] = 8'h00;
mem[16'hC37B] = 8'h00;
mem[16'hC37C] = 8'h00;
mem[16'hC37D] = 8'h00;
mem[16'hC37E] = 8'h00;
mem[16'hC37F] = 8'h00;
mem[16'hC380] = 8'h00;
mem[16'hC381] = 8'h00;
mem[16'hC382] = 8'h00;
mem[16'hC383] = 8'h00;
mem[16'hC384] = 8'h00;
mem[16'hC385] = 8'h00;
mem[16'hC386] = 8'h00;
mem[16'hC387] = 8'h00;
mem[16'hC388] = 8'h00;
mem[16'hC389] = 8'h00;
mem[16'hC38A] = 8'h00;
mem[16'hC38B] = 8'h00;
mem[16'hC38C] = 8'h00;
mem[16'hC38D] = 8'h00;
mem[16'hC38E] = 8'h00;
mem[16'hC38F] = 8'h00;
mem[16'hC390] = 8'h00;
mem[16'hC391] = 8'h00;
mem[16'hC392] = 8'h00;
mem[16'hC393] = 8'h00;
mem[16'hC394] = 8'h00;
mem[16'hC395] = 8'h00;
mem[16'hC396] = 8'h00;
mem[16'hC397] = 8'h00;
mem[16'hC398] = 8'h00;
mem[16'hC399] = 8'h00;
mem[16'hC39A] = 8'h00;
mem[16'hC39B] = 8'h00;
mem[16'hC39C] = 8'h00;
mem[16'hC39D] = 8'h00;
mem[16'hC39E] = 8'h00;
mem[16'hC39F] = 8'h00;
mem[16'hC3A0] = 8'h00;
mem[16'hC3A1] = 8'h00;
mem[16'hC3A2] = 8'h00;
mem[16'hC3A3] = 8'h00;
mem[16'hC3A4] = 8'h00;
mem[16'hC3A5] = 8'h00;
mem[16'hC3A6] = 8'h00;
mem[16'hC3A7] = 8'h00;
mem[16'hC3A8] = 8'h00;
mem[16'hC3A9] = 8'h00;
mem[16'hC3AA] = 8'h00;
mem[16'hC3AB] = 8'h00;
mem[16'hC3AC] = 8'h00;
mem[16'hC3AD] = 8'h00;
mem[16'hC3AE] = 8'h00;
mem[16'hC3AF] = 8'h00;
mem[16'hC3B0] = 8'h00;
mem[16'hC3B1] = 8'h00;
mem[16'hC3B2] = 8'h00;
mem[16'hC3B3] = 8'h00;
mem[16'hC3B4] = 8'h00;
mem[16'hC3B5] = 8'h00;
mem[16'hC3B6] = 8'h00;
mem[16'hC3B7] = 8'h00;
mem[16'hC3B8] = 8'h00;
mem[16'hC3B9] = 8'h00;
mem[16'hC3BA] = 8'h00;
mem[16'hC3BB] = 8'h00;
mem[16'hC3BC] = 8'h00;
mem[16'hC3BD] = 8'h00;
mem[16'hC3BE] = 8'h00;
mem[16'hC3BF] = 8'h00;
mem[16'hC3C0] = 8'h00;
mem[16'hC3C1] = 8'h00;
mem[16'hC3C2] = 8'h00;
mem[16'hC3C3] = 8'h00;
mem[16'hC3C4] = 8'h00;
mem[16'hC3C5] = 8'h00;
mem[16'hC3C6] = 8'h00;
mem[16'hC3C7] = 8'h00;
mem[16'hC3C8] = 8'h00;
mem[16'hC3C9] = 8'h00;
mem[16'hC3CA] = 8'h00;
mem[16'hC3CB] = 8'h00;
mem[16'hC3CC] = 8'h00;
mem[16'hC3CD] = 8'h00;
mem[16'hC3CE] = 8'h00;
mem[16'hC3CF] = 8'h00;
mem[16'hC3D0] = 8'h00;
mem[16'hC3D1] = 8'h00;
mem[16'hC3D2] = 8'h00;
mem[16'hC3D3] = 8'h00;
mem[16'hC3D4] = 8'h00;
mem[16'hC3D5] = 8'h00;
mem[16'hC3D6] = 8'h00;
mem[16'hC3D7] = 8'h00;
mem[16'hC3D8] = 8'h00;
mem[16'hC3D9] = 8'h00;
mem[16'hC3DA] = 8'h00;
mem[16'hC3DB] = 8'h00;
mem[16'hC3DC] = 8'h00;
mem[16'hC3DD] = 8'h00;
mem[16'hC3DE] = 8'h00;
mem[16'hC3DF] = 8'h00;
mem[16'hC3E0] = 8'h00;
mem[16'hC3E1] = 8'h00;
mem[16'hC3E2] = 8'h00;
mem[16'hC3E3] = 8'h00;
mem[16'hC3E4] = 8'h00;
mem[16'hC3E5] = 8'h00;
mem[16'hC3E6] = 8'h00;
mem[16'hC3E7] = 8'h00;
mem[16'hC3E8] = 8'h00;
mem[16'hC3E9] = 8'h00;
mem[16'hC3EA] = 8'h00;
mem[16'hC3EB] = 8'h00;
mem[16'hC3EC] = 8'h00;
mem[16'hC3ED] = 8'h00;
mem[16'hC3EE] = 8'h00;
mem[16'hC3EF] = 8'h00;
mem[16'hC3F0] = 8'h00;
mem[16'hC3F1] = 8'h00;
mem[16'hC3F2] = 8'h00;
mem[16'hC3F3] = 8'h00;
mem[16'hC3F4] = 8'h00;
mem[16'hC3F5] = 8'h00;
mem[16'hC3F6] = 8'h00;
mem[16'hC3F7] = 8'h00;
mem[16'hC3F8] = 8'h00;
mem[16'hC3F9] = 8'h00;
mem[16'hC3FA] = 8'h00;
mem[16'hC3FB] = 8'h00;
mem[16'hC3FC] = 8'h00;
mem[16'hC3FD] = 8'h00;
mem[16'hC3FE] = 8'h00;
mem[16'hC3FF] = 8'h00;
mem[16'hC400] = 8'h00;
mem[16'hC401] = 8'h00;
mem[16'hC402] = 8'h00;
mem[16'hC403] = 8'h00;
mem[16'hC404] = 8'h00;
mem[16'hC405] = 8'h00;
mem[16'hC406] = 8'h00;
mem[16'hC407] = 8'h00;
mem[16'hC408] = 8'h00;
mem[16'hC409] = 8'h00;
mem[16'hC40A] = 8'h00;
mem[16'hC40B] = 8'h00;
mem[16'hC40C] = 8'h00;
mem[16'hC40D] = 8'h00;
mem[16'hC40E] = 8'h00;
mem[16'hC40F] = 8'h00;
mem[16'hC410] = 8'h00;
mem[16'hC411] = 8'h00;
mem[16'hC412] = 8'h00;
mem[16'hC413] = 8'h00;
mem[16'hC414] = 8'h00;
mem[16'hC415] = 8'h00;
mem[16'hC416] = 8'h00;
mem[16'hC417] = 8'h00;
mem[16'hC418] = 8'h00;
mem[16'hC419] = 8'h00;
mem[16'hC41A] = 8'h00;
mem[16'hC41B] = 8'h00;
mem[16'hC41C] = 8'h00;
mem[16'hC41D] = 8'h00;
mem[16'hC41E] = 8'h00;
mem[16'hC41F] = 8'h00;
mem[16'hC420] = 8'h00;
mem[16'hC421] = 8'h00;
mem[16'hC422] = 8'h00;
mem[16'hC423] = 8'h00;
mem[16'hC424] = 8'h00;
mem[16'hC425] = 8'h00;
mem[16'hC426] = 8'h00;
mem[16'hC427] = 8'h00;
mem[16'hC428] = 8'h00;
mem[16'hC429] = 8'h00;
mem[16'hC42A] = 8'h00;
mem[16'hC42B] = 8'h00;
mem[16'hC42C] = 8'h00;
mem[16'hC42D] = 8'h00;
mem[16'hC42E] = 8'h00;
mem[16'hC42F] = 8'h00;
mem[16'hC430] = 8'h00;
mem[16'hC431] = 8'h00;
mem[16'hC432] = 8'h00;
mem[16'hC433] = 8'h00;
mem[16'hC434] = 8'h00;
mem[16'hC435] = 8'h00;
mem[16'hC436] = 8'h00;
mem[16'hC437] = 8'h00;
mem[16'hC438] = 8'h00;
mem[16'hC439] = 8'h00;
mem[16'hC43A] = 8'h00;
mem[16'hC43B] = 8'h00;
mem[16'hC43C] = 8'h00;
mem[16'hC43D] = 8'h00;
mem[16'hC43E] = 8'h00;
mem[16'hC43F] = 8'h00;
mem[16'hC440] = 8'h00;
mem[16'hC441] = 8'h00;
mem[16'hC442] = 8'h00;
mem[16'hC443] = 8'h00;
mem[16'hC444] = 8'h00;
mem[16'hC445] = 8'h00;
mem[16'hC446] = 8'h00;
mem[16'hC447] = 8'h00;
mem[16'hC448] = 8'h00;
mem[16'hC449] = 8'h00;
mem[16'hC44A] = 8'h00;
mem[16'hC44B] = 8'h00;
mem[16'hC44C] = 8'h00;
mem[16'hC44D] = 8'h00;
mem[16'hC44E] = 8'h00;
mem[16'hC44F] = 8'h00;
mem[16'hC450] = 8'h00;
mem[16'hC451] = 8'h00;
mem[16'hC452] = 8'h00;
mem[16'hC453] = 8'h00;
mem[16'hC454] = 8'h00;
mem[16'hC455] = 8'h00;
mem[16'hC456] = 8'h00;
mem[16'hC457] = 8'h00;
mem[16'hC458] = 8'h00;
mem[16'hC459] = 8'h00;
mem[16'hC45A] = 8'h00;
mem[16'hC45B] = 8'h00;
mem[16'hC45C] = 8'h00;
mem[16'hC45D] = 8'h00;
mem[16'hC45E] = 8'h00;
mem[16'hC45F] = 8'h00;
mem[16'hC460] = 8'h00;
mem[16'hC461] = 8'h00;
mem[16'hC462] = 8'h00;
mem[16'hC463] = 8'h00;
mem[16'hC464] = 8'h00;
mem[16'hC465] = 8'h00;
mem[16'hC466] = 8'h00;
mem[16'hC467] = 8'h00;
mem[16'hC468] = 8'h00;
mem[16'hC469] = 8'h00;
mem[16'hC46A] = 8'h00;
mem[16'hC46B] = 8'h00;
mem[16'hC46C] = 8'h00;
mem[16'hC46D] = 8'h00;
mem[16'hC46E] = 8'h00;
mem[16'hC46F] = 8'h00;
mem[16'hC470] = 8'h00;
mem[16'hC471] = 8'h00;
mem[16'hC472] = 8'h00;
mem[16'hC473] = 8'h00;
mem[16'hC474] = 8'h00;
mem[16'hC475] = 8'h00;
mem[16'hC476] = 8'h00;
mem[16'hC477] = 8'h00;
mem[16'hC478] = 8'h00;
mem[16'hC479] = 8'h00;
mem[16'hC47A] = 8'h00;
mem[16'hC47B] = 8'h00;
mem[16'hC47C] = 8'h00;
mem[16'hC47D] = 8'h00;
mem[16'hC47E] = 8'h00;
mem[16'hC47F] = 8'h00;
mem[16'hC480] = 8'h00;
mem[16'hC481] = 8'h00;
mem[16'hC482] = 8'h00;
mem[16'hC483] = 8'h00;
mem[16'hC484] = 8'h00;
mem[16'hC485] = 8'h00;
mem[16'hC486] = 8'h00;
mem[16'hC487] = 8'h00;
mem[16'hC488] = 8'h00;
mem[16'hC489] = 8'h00;
mem[16'hC48A] = 8'h00;
mem[16'hC48B] = 8'h00;
mem[16'hC48C] = 8'h00;
mem[16'hC48D] = 8'h00;
mem[16'hC48E] = 8'h00;
mem[16'hC48F] = 8'h00;
mem[16'hC490] = 8'h00;
mem[16'hC491] = 8'h00;
mem[16'hC492] = 8'h00;
mem[16'hC493] = 8'h00;
mem[16'hC494] = 8'h00;
mem[16'hC495] = 8'h00;
mem[16'hC496] = 8'h00;
mem[16'hC497] = 8'h00;
mem[16'hC498] = 8'h00;
mem[16'hC499] = 8'h00;
mem[16'hC49A] = 8'h00;
mem[16'hC49B] = 8'h00;
mem[16'hC49C] = 8'h00;
mem[16'hC49D] = 8'h00;
mem[16'hC49E] = 8'h00;
mem[16'hC49F] = 8'h00;
mem[16'hC4A0] = 8'h00;
mem[16'hC4A1] = 8'h00;
mem[16'hC4A2] = 8'h00;
mem[16'hC4A3] = 8'h00;
mem[16'hC4A4] = 8'h00;
mem[16'hC4A5] = 8'h00;
mem[16'hC4A6] = 8'h00;
mem[16'hC4A7] = 8'h00;
mem[16'hC4A8] = 8'h00;
mem[16'hC4A9] = 8'h00;
mem[16'hC4AA] = 8'h00;
mem[16'hC4AB] = 8'h00;
mem[16'hC4AC] = 8'h00;
mem[16'hC4AD] = 8'h00;
mem[16'hC4AE] = 8'h00;
mem[16'hC4AF] = 8'h00;
mem[16'hC4B0] = 8'h00;
mem[16'hC4B1] = 8'h00;
mem[16'hC4B2] = 8'h00;
mem[16'hC4B3] = 8'h00;
mem[16'hC4B4] = 8'h00;
mem[16'hC4B5] = 8'h00;
mem[16'hC4B6] = 8'h00;
mem[16'hC4B7] = 8'h00;
mem[16'hC4B8] = 8'h00;
mem[16'hC4B9] = 8'h00;
mem[16'hC4BA] = 8'h00;
mem[16'hC4BB] = 8'h00;
mem[16'hC4BC] = 8'h00;
mem[16'hC4BD] = 8'h00;
mem[16'hC4BE] = 8'h00;
mem[16'hC4BF] = 8'h00;
mem[16'hC4C0] = 8'h00;
mem[16'hC4C1] = 8'h00;
mem[16'hC4C2] = 8'h00;
mem[16'hC4C3] = 8'h00;
mem[16'hC4C4] = 8'h00;
mem[16'hC4C5] = 8'h00;
mem[16'hC4C6] = 8'h00;
mem[16'hC4C7] = 8'h00;
mem[16'hC4C8] = 8'h00;
mem[16'hC4C9] = 8'h00;
mem[16'hC4CA] = 8'h00;
mem[16'hC4CB] = 8'h00;
mem[16'hC4CC] = 8'h00;
mem[16'hC4CD] = 8'h00;
mem[16'hC4CE] = 8'h00;
mem[16'hC4CF] = 8'h00;
mem[16'hC4D0] = 8'h00;
mem[16'hC4D1] = 8'h00;
mem[16'hC4D2] = 8'h00;
mem[16'hC4D3] = 8'h00;
mem[16'hC4D4] = 8'h00;
mem[16'hC4D5] = 8'h00;
mem[16'hC4D6] = 8'h00;
mem[16'hC4D7] = 8'h00;
mem[16'hC4D8] = 8'h00;
mem[16'hC4D9] = 8'h00;
mem[16'hC4DA] = 8'h00;
mem[16'hC4DB] = 8'h00;
mem[16'hC4DC] = 8'h00;
mem[16'hC4DD] = 8'h00;
mem[16'hC4DE] = 8'h00;
mem[16'hC4DF] = 8'h00;
mem[16'hC4E0] = 8'h00;
mem[16'hC4E1] = 8'h00;
mem[16'hC4E2] = 8'h00;
mem[16'hC4E3] = 8'h00;
mem[16'hC4E4] = 8'h00;
mem[16'hC4E5] = 8'h00;
mem[16'hC4E6] = 8'h00;
mem[16'hC4E7] = 8'h00;
mem[16'hC4E8] = 8'h00;
mem[16'hC4E9] = 8'h00;
mem[16'hC4EA] = 8'h00;
mem[16'hC4EB] = 8'h00;
mem[16'hC4EC] = 8'h00;
mem[16'hC4ED] = 8'h00;
mem[16'hC4EE] = 8'h00;
mem[16'hC4EF] = 8'h00;
mem[16'hC4F0] = 8'h00;
mem[16'hC4F1] = 8'h00;
mem[16'hC4F2] = 8'h00;
mem[16'hC4F3] = 8'h00;
mem[16'hC4F4] = 8'h00;
mem[16'hC4F5] = 8'h00;
mem[16'hC4F6] = 8'h00;
mem[16'hC4F7] = 8'h00;
mem[16'hC4F8] = 8'h00;
mem[16'hC4F9] = 8'h00;
mem[16'hC4FA] = 8'h00;
mem[16'hC4FB] = 8'h00;
mem[16'hC4FC] = 8'h00;
mem[16'hC4FD] = 8'h00;
mem[16'hC4FE] = 8'h00;
mem[16'hC4FF] = 8'h00;
mem[16'hC500] = 8'h00;
mem[16'hC501] = 8'h00;
mem[16'hC502] = 8'h00;
mem[16'hC503] = 8'h00;
mem[16'hC504] = 8'h00;
mem[16'hC505] = 8'h00;
mem[16'hC506] = 8'h00;
mem[16'hC507] = 8'h00;
mem[16'hC508] = 8'h00;
mem[16'hC509] = 8'h00;
mem[16'hC50A] = 8'h00;
mem[16'hC50B] = 8'h00;
mem[16'hC50C] = 8'h00;
mem[16'hC50D] = 8'h00;
mem[16'hC50E] = 8'h00;
mem[16'hC50F] = 8'h00;
mem[16'hC510] = 8'h00;
mem[16'hC511] = 8'h00;
mem[16'hC512] = 8'h00;
mem[16'hC513] = 8'h00;
mem[16'hC514] = 8'h00;
mem[16'hC515] = 8'h00;
mem[16'hC516] = 8'h00;
mem[16'hC517] = 8'h00;
mem[16'hC518] = 8'h00;
mem[16'hC519] = 8'h00;
mem[16'hC51A] = 8'h00;
mem[16'hC51B] = 8'h00;
mem[16'hC51C] = 8'h00;
mem[16'hC51D] = 8'h00;
mem[16'hC51E] = 8'h00;
mem[16'hC51F] = 8'h00;
mem[16'hC520] = 8'h00;
mem[16'hC521] = 8'h00;
mem[16'hC522] = 8'h00;
mem[16'hC523] = 8'h00;
mem[16'hC524] = 8'h00;
mem[16'hC525] = 8'h00;
mem[16'hC526] = 8'h00;
mem[16'hC527] = 8'h00;
mem[16'hC528] = 8'h00;
mem[16'hC529] = 8'h00;
mem[16'hC52A] = 8'h00;
mem[16'hC52B] = 8'h00;
mem[16'hC52C] = 8'h00;
mem[16'hC52D] = 8'h00;
mem[16'hC52E] = 8'h00;
mem[16'hC52F] = 8'h00;
mem[16'hC530] = 8'h00;
mem[16'hC531] = 8'h00;
mem[16'hC532] = 8'h00;
mem[16'hC533] = 8'h00;
mem[16'hC534] = 8'h00;
mem[16'hC535] = 8'h00;
mem[16'hC536] = 8'h00;
mem[16'hC537] = 8'h00;
mem[16'hC538] = 8'h00;
mem[16'hC539] = 8'h00;
mem[16'hC53A] = 8'h00;
mem[16'hC53B] = 8'h00;
mem[16'hC53C] = 8'h00;
mem[16'hC53D] = 8'h00;
mem[16'hC53E] = 8'h00;
mem[16'hC53F] = 8'h00;
mem[16'hC540] = 8'h00;
mem[16'hC541] = 8'h00;
mem[16'hC542] = 8'h00;
mem[16'hC543] = 8'h00;
mem[16'hC544] = 8'h00;
mem[16'hC545] = 8'h00;
mem[16'hC546] = 8'h00;
mem[16'hC547] = 8'h00;
mem[16'hC548] = 8'h00;
mem[16'hC549] = 8'h00;
mem[16'hC54A] = 8'h00;
mem[16'hC54B] = 8'h00;
mem[16'hC54C] = 8'h00;
mem[16'hC54D] = 8'h00;
mem[16'hC54E] = 8'h00;
mem[16'hC54F] = 8'h00;
mem[16'hC550] = 8'h00;
mem[16'hC551] = 8'h00;
mem[16'hC552] = 8'h00;
mem[16'hC553] = 8'h00;
mem[16'hC554] = 8'h00;
mem[16'hC555] = 8'h00;
mem[16'hC556] = 8'h00;
mem[16'hC557] = 8'h00;
mem[16'hC558] = 8'h00;
mem[16'hC559] = 8'h00;
mem[16'hC55A] = 8'h00;
mem[16'hC55B] = 8'h00;
mem[16'hC55C] = 8'h00;
mem[16'hC55D] = 8'h00;
mem[16'hC55E] = 8'h00;
mem[16'hC55F] = 8'h00;
mem[16'hC560] = 8'h00;
mem[16'hC561] = 8'h00;
mem[16'hC562] = 8'h00;
mem[16'hC563] = 8'h00;
mem[16'hC564] = 8'h00;
mem[16'hC565] = 8'h00;
mem[16'hC566] = 8'h00;
mem[16'hC567] = 8'h00;
mem[16'hC568] = 8'h00;
mem[16'hC569] = 8'h00;
mem[16'hC56A] = 8'h00;
mem[16'hC56B] = 8'h00;
mem[16'hC56C] = 8'h00;
mem[16'hC56D] = 8'h00;
mem[16'hC56E] = 8'h00;
mem[16'hC56F] = 8'h00;
mem[16'hC570] = 8'h00;
mem[16'hC571] = 8'h00;
mem[16'hC572] = 8'h00;
mem[16'hC573] = 8'h00;
mem[16'hC574] = 8'h00;
mem[16'hC575] = 8'h00;
mem[16'hC576] = 8'h00;
mem[16'hC577] = 8'h00;
mem[16'hC578] = 8'h00;
mem[16'hC579] = 8'h00;
mem[16'hC57A] = 8'h00;
mem[16'hC57B] = 8'h00;
mem[16'hC57C] = 8'h00;
mem[16'hC57D] = 8'h00;
mem[16'hC57E] = 8'h00;
mem[16'hC57F] = 8'h00;
mem[16'hC580] = 8'h00;
mem[16'hC581] = 8'h00;
mem[16'hC582] = 8'h00;
mem[16'hC583] = 8'h00;
mem[16'hC584] = 8'h00;
mem[16'hC585] = 8'h00;
mem[16'hC586] = 8'h00;
mem[16'hC587] = 8'h00;
mem[16'hC588] = 8'h00;
mem[16'hC589] = 8'h00;
mem[16'hC58A] = 8'h00;
mem[16'hC58B] = 8'h00;
mem[16'hC58C] = 8'h00;
mem[16'hC58D] = 8'h00;
mem[16'hC58E] = 8'h00;
mem[16'hC58F] = 8'h00;
mem[16'hC590] = 8'h00;
mem[16'hC591] = 8'h00;
mem[16'hC592] = 8'h00;
mem[16'hC593] = 8'h00;
mem[16'hC594] = 8'h00;
mem[16'hC595] = 8'h00;
mem[16'hC596] = 8'h00;
mem[16'hC597] = 8'h00;
mem[16'hC598] = 8'h00;
mem[16'hC599] = 8'h00;
mem[16'hC59A] = 8'h00;
mem[16'hC59B] = 8'h00;
mem[16'hC59C] = 8'h00;
mem[16'hC59D] = 8'h00;
mem[16'hC59E] = 8'h00;
mem[16'hC59F] = 8'h00;
mem[16'hC5A0] = 8'h00;
mem[16'hC5A1] = 8'h00;
mem[16'hC5A2] = 8'h00;
mem[16'hC5A3] = 8'h00;
mem[16'hC5A4] = 8'h00;
mem[16'hC5A5] = 8'h00;
mem[16'hC5A6] = 8'h00;
mem[16'hC5A7] = 8'h00;
mem[16'hC5A8] = 8'h00;
mem[16'hC5A9] = 8'h00;
mem[16'hC5AA] = 8'h00;
mem[16'hC5AB] = 8'h00;
mem[16'hC5AC] = 8'h00;
mem[16'hC5AD] = 8'h00;
mem[16'hC5AE] = 8'h00;
mem[16'hC5AF] = 8'h00;
mem[16'hC5B0] = 8'h00;
mem[16'hC5B1] = 8'h00;
mem[16'hC5B2] = 8'h00;
mem[16'hC5B3] = 8'h00;
mem[16'hC5B4] = 8'h00;
mem[16'hC5B5] = 8'h00;
mem[16'hC5B6] = 8'h00;
mem[16'hC5B7] = 8'h00;
mem[16'hC5B8] = 8'h00;
mem[16'hC5B9] = 8'h00;
mem[16'hC5BA] = 8'h00;
mem[16'hC5BB] = 8'h00;
mem[16'hC5BC] = 8'h00;
mem[16'hC5BD] = 8'h00;
mem[16'hC5BE] = 8'h00;
mem[16'hC5BF] = 8'h00;
mem[16'hC5C0] = 8'h00;
mem[16'hC5C1] = 8'h00;
mem[16'hC5C2] = 8'h00;
mem[16'hC5C3] = 8'h00;
mem[16'hC5C4] = 8'h00;
mem[16'hC5C5] = 8'h00;
mem[16'hC5C6] = 8'h00;
mem[16'hC5C7] = 8'h00;
mem[16'hC5C8] = 8'h00;
mem[16'hC5C9] = 8'h00;
mem[16'hC5CA] = 8'h00;
mem[16'hC5CB] = 8'h00;
mem[16'hC5CC] = 8'h00;
mem[16'hC5CD] = 8'h00;
mem[16'hC5CE] = 8'h00;
mem[16'hC5CF] = 8'h00;
mem[16'hC5D0] = 8'h00;
mem[16'hC5D1] = 8'h00;
mem[16'hC5D2] = 8'h00;
mem[16'hC5D3] = 8'h00;
mem[16'hC5D4] = 8'h00;
mem[16'hC5D5] = 8'h00;
mem[16'hC5D6] = 8'h00;
mem[16'hC5D7] = 8'h00;
mem[16'hC5D8] = 8'h00;
mem[16'hC5D9] = 8'h00;
mem[16'hC5DA] = 8'h00;
mem[16'hC5DB] = 8'h00;
mem[16'hC5DC] = 8'h00;
mem[16'hC5DD] = 8'h00;
mem[16'hC5DE] = 8'h00;
mem[16'hC5DF] = 8'h00;
mem[16'hC5E0] = 8'h00;
mem[16'hC5E1] = 8'h00;
mem[16'hC5E2] = 8'h00;
mem[16'hC5E3] = 8'h00;
mem[16'hC5E4] = 8'h00;
mem[16'hC5E5] = 8'h00;
mem[16'hC5E6] = 8'h00;
mem[16'hC5E7] = 8'h00;
mem[16'hC5E8] = 8'h00;
mem[16'hC5E9] = 8'h00;
mem[16'hC5EA] = 8'h00;
mem[16'hC5EB] = 8'h00;
mem[16'hC5EC] = 8'h00;
mem[16'hC5ED] = 8'h00;
mem[16'hC5EE] = 8'h00;
mem[16'hC5EF] = 8'h00;
mem[16'hC5F0] = 8'h00;
mem[16'hC5F1] = 8'h00;
mem[16'hC5F2] = 8'h00;
mem[16'hC5F3] = 8'h00;
mem[16'hC5F4] = 8'h00;
mem[16'hC5F5] = 8'h00;
mem[16'hC5F6] = 8'h00;
mem[16'hC5F7] = 8'h00;
mem[16'hC5F8] = 8'h00;
mem[16'hC5F9] = 8'h00;
mem[16'hC5FA] = 8'h00;
mem[16'hC5FB] = 8'h00;
mem[16'hC5FC] = 8'h00;
mem[16'hC5FD] = 8'h00;
mem[16'hC5FE] = 8'h00;
mem[16'hC5FF] = 8'h00;
mem[16'hC600] = 8'hA2;
mem[16'hC601] = 8'h20;
mem[16'hC602] = 8'hA0;
mem[16'hC603] = 8'h00;
mem[16'hC604] = 8'hA2;
mem[16'hC605] = 8'h03;
mem[16'hC606] = 8'h86;
mem[16'hC607] = 8'h3C;
mem[16'hC608] = 8'h8A;
mem[16'hC609] = 8'h0A;
mem[16'hC60A] = 8'h24;
mem[16'hC60B] = 8'h3C;
mem[16'hC60C] = 8'hF0;
mem[16'hC60D] = 8'h10;
mem[16'hC60E] = 8'h05;
mem[16'hC60F] = 8'h3C;
mem[16'hC610] = 8'h49;
mem[16'hC611] = 8'hFF;
mem[16'hC612] = 8'h29;
mem[16'hC613] = 8'h7E;
mem[16'hC614] = 8'hB0;
mem[16'hC615] = 8'h08;
mem[16'hC616] = 8'h4A;
mem[16'hC617] = 8'hD0;
mem[16'hC618] = 8'hFB;
mem[16'hC619] = 8'h98;
mem[16'hC61A] = 8'h9D;
mem[16'hC61B] = 8'h56;
mem[16'hC61C] = 8'h03;
mem[16'hC61D] = 8'hC8;
mem[16'hC61E] = 8'hE8;
mem[16'hC61F] = 8'h10;
mem[16'hC620] = 8'hE5;
mem[16'hC621] = 8'h20;
mem[16'hC622] = 8'h58;
mem[16'hC623] = 8'hFF;
mem[16'hC624] = 8'hBA;
mem[16'hC625] = 8'hBD;
mem[16'hC626] = 8'h00;
mem[16'hC627] = 8'h01;
mem[16'hC628] = 8'h0A;
mem[16'hC629] = 8'h0A;
mem[16'hC62A] = 8'h0A;
mem[16'hC62B] = 8'h0A;
mem[16'hC62C] = 8'h85;
mem[16'hC62D] = 8'h2B;
mem[16'hC62E] = 8'hAA;
mem[16'hC62F] = 8'hBD;
mem[16'hC630] = 8'h8E;
mem[16'hC631] = 8'hC0;
mem[16'hC632] = 8'hBD;
mem[16'hC633] = 8'h8C;
mem[16'hC634] = 8'hC0;
mem[16'hC635] = 8'hBD;
mem[16'hC636] = 8'h8A;
mem[16'hC637] = 8'hC0;
mem[16'hC638] = 8'hBD;
mem[16'hC639] = 8'h89;
mem[16'hC63A] = 8'hC0;
mem[16'hC63B] = 8'hA0;
mem[16'hC63C] = 8'h50;
mem[16'hC63D] = 8'hBD;
mem[16'hC63E] = 8'h80;
mem[16'hC63F] = 8'hC0;
mem[16'hC640] = 8'h98;
mem[16'hC641] = 8'h29;
mem[16'hC642] = 8'h03;
mem[16'hC643] = 8'h0A;
mem[16'hC644] = 8'h05;
mem[16'hC645] = 8'h2B;
mem[16'hC646] = 8'hAA;
mem[16'hC647] = 8'hBD;
mem[16'hC648] = 8'h81;
mem[16'hC649] = 8'hC0;
mem[16'hC64A] = 8'hA9;
mem[16'hC64B] = 8'h56;
mem[16'hC64C] = 8'h20;
mem[16'hC64D] = 8'hA8;
mem[16'hC64E] = 8'hFC;
mem[16'hC64F] = 8'h88;
mem[16'hC650] = 8'h10;
mem[16'hC651] = 8'hEB;
mem[16'hC652] = 8'h85;
mem[16'hC653] = 8'h26;
mem[16'hC654] = 8'h85;
mem[16'hC655] = 8'h3D;
mem[16'hC656] = 8'h85;
mem[16'hC657] = 8'h41;
mem[16'hC658] = 8'hA9;
mem[16'hC659] = 8'h08;
mem[16'hC65A] = 8'h85;
mem[16'hC65B] = 8'h27;
mem[16'hC65C] = 8'h18;
mem[16'hC65D] = 8'h08;
mem[16'hC65E] = 8'hBD;
mem[16'hC65F] = 8'h8C;
mem[16'hC660] = 8'hC0;
mem[16'hC661] = 8'h10;
mem[16'hC662] = 8'hFB;
mem[16'hC663] = 8'h49;
mem[16'hC664] = 8'hD5;
mem[16'hC665] = 8'hD0;
mem[16'hC666] = 8'hF7;
mem[16'hC667] = 8'hBD;
mem[16'hC668] = 8'h8C;
mem[16'hC669] = 8'hC0;
mem[16'hC66A] = 8'h10;
mem[16'hC66B] = 8'hFB;
mem[16'hC66C] = 8'hC9;
mem[16'hC66D] = 8'hAA;
mem[16'hC66E] = 8'hD0;
mem[16'hC66F] = 8'hF3;
mem[16'hC670] = 8'hEA;
mem[16'hC671] = 8'hBD;
mem[16'hC672] = 8'h8C;
mem[16'hC673] = 8'hC0;
mem[16'hC674] = 8'h10;
mem[16'hC675] = 8'hFB;
mem[16'hC676] = 8'hC9;
mem[16'hC677] = 8'h96;
mem[16'hC678] = 8'hF0;
mem[16'hC679] = 8'h09;
mem[16'hC67A] = 8'h28;
mem[16'hC67B] = 8'h90;
mem[16'hC67C] = 8'hDF;
mem[16'hC67D] = 8'h49;
mem[16'hC67E] = 8'hAD;
mem[16'hC67F] = 8'hF0;
mem[16'hC680] = 8'h25;
mem[16'hC681] = 8'hD0;
mem[16'hC682] = 8'hD9;
mem[16'hC683] = 8'hA0;
mem[16'hC684] = 8'h03;
mem[16'hC685] = 8'h85;
mem[16'hC686] = 8'h40;
mem[16'hC687] = 8'hBD;
mem[16'hC688] = 8'h8C;
mem[16'hC689] = 8'hC0;
mem[16'hC68A] = 8'h10;
mem[16'hC68B] = 8'hFB;
mem[16'hC68C] = 8'h2A;
mem[16'hC68D] = 8'h85;
mem[16'hC68E] = 8'h3C;
mem[16'hC68F] = 8'hBD;
mem[16'hC690] = 8'h8C;
mem[16'hC691] = 8'hC0;
mem[16'hC692] = 8'h10;
mem[16'hC693] = 8'hFB;
mem[16'hC694] = 8'h25;
mem[16'hC695] = 8'h3C;
mem[16'hC696] = 8'h88;
mem[16'hC697] = 8'hD0;
mem[16'hC698] = 8'hEC;
mem[16'hC699] = 8'h28;
mem[16'hC69A] = 8'hC5;
mem[16'hC69B] = 8'h3D;
mem[16'hC69C] = 8'hD0;
mem[16'hC69D] = 8'hBE;
mem[16'hC69E] = 8'hA5;
mem[16'hC69F] = 8'h40;
mem[16'hC6A0] = 8'hC5;
mem[16'hC6A1] = 8'h41;
mem[16'hC6A2] = 8'hD0;
mem[16'hC6A3] = 8'hB8;
mem[16'hC6A4] = 8'hB0;
mem[16'hC6A5] = 8'hB7;
mem[16'hC6A6] = 8'hA0;
mem[16'hC6A7] = 8'h56;
mem[16'hC6A8] = 8'h84;
mem[16'hC6A9] = 8'h3C;
mem[16'hC6AA] = 8'hBC;
mem[16'hC6AB] = 8'h8C;
mem[16'hC6AC] = 8'hC0;
mem[16'hC6AD] = 8'h10;
mem[16'hC6AE] = 8'hFB;
mem[16'hC6AF] = 8'h59;
mem[16'hC6B0] = 8'hD6;
mem[16'hC6B1] = 8'h02;
mem[16'hC6B2] = 8'hA4;
mem[16'hC6B3] = 8'h3C;
mem[16'hC6B4] = 8'h88;
mem[16'hC6B5] = 8'h99;
mem[16'hC6B6] = 8'h00;
mem[16'hC6B7] = 8'h03;
mem[16'hC6B8] = 8'hD0;
mem[16'hC6B9] = 8'hEE;
mem[16'hC6BA] = 8'h84;
mem[16'hC6BB] = 8'h3C;
mem[16'hC6BC] = 8'hBC;
mem[16'hC6BD] = 8'h8C;
mem[16'hC6BE] = 8'hC0;
mem[16'hC6BF] = 8'h10;
mem[16'hC6C0] = 8'hFB;
mem[16'hC6C1] = 8'h59;
mem[16'hC6C2] = 8'hD6;
mem[16'hC6C3] = 8'h02;
mem[16'hC6C4] = 8'hA4;
mem[16'hC6C5] = 8'h3C;
mem[16'hC6C6] = 8'h91;
mem[16'hC6C7] = 8'h26;
mem[16'hC6C8] = 8'hC8;
mem[16'hC6C9] = 8'hD0;
mem[16'hC6CA] = 8'hEF;
mem[16'hC6CB] = 8'hBC;
mem[16'hC6CC] = 8'h8C;
mem[16'hC6CD] = 8'hC0;
mem[16'hC6CE] = 8'h10;
mem[16'hC6CF] = 8'hFB;
mem[16'hC6D0] = 8'h59;
mem[16'hC6D1] = 8'hD6;
mem[16'hC6D2] = 8'h02;
mem[16'hC6D3] = 8'hD0;
mem[16'hC6D4] = 8'h87;
mem[16'hC6D5] = 8'hA0;
mem[16'hC6D6] = 8'h00;
mem[16'hC6D7] = 8'hA2;
mem[16'hC6D8] = 8'h56;
mem[16'hC6D9] = 8'hCA;
mem[16'hC6DA] = 8'h30;
mem[16'hC6DB] = 8'hFB;
mem[16'hC6DC] = 8'hB1;
mem[16'hC6DD] = 8'h26;
mem[16'hC6DE] = 8'h5E;
mem[16'hC6DF] = 8'h00;
mem[16'hC6E0] = 8'h03;
mem[16'hC6E1] = 8'h2A;
mem[16'hC6E2] = 8'h5E;
mem[16'hC6E3] = 8'h00;
mem[16'hC6E4] = 8'h03;
mem[16'hC6E5] = 8'h2A;
mem[16'hC6E6] = 8'h91;
mem[16'hC6E7] = 8'h26;
mem[16'hC6E8] = 8'hC8;
mem[16'hC6E9] = 8'hD0;
mem[16'hC6EA] = 8'hEE;
mem[16'hC6EB] = 8'hE6;
mem[16'hC6EC] = 8'h27;
mem[16'hC6ED] = 8'hE6;
mem[16'hC6EE] = 8'h3D;
mem[16'hC6EF] = 8'hA5;
mem[16'hC6F0] = 8'h3D;
mem[16'hC6F1] = 8'hCD;
mem[16'hC6F2] = 8'h00;
mem[16'hC6F3] = 8'h08;
mem[16'hC6F4] = 8'hA6;
mem[16'hC6F5] = 8'h2B;
mem[16'hC6F6] = 8'h90;
mem[16'hC6F7] = 8'hDB;
mem[16'hC6F8] = 8'h4C;
mem[16'hC6F9] = 8'h01;
mem[16'hC6FA] = 8'h08;
mem[16'hC6FB] = 8'h00;
mem[16'hC6FC] = 8'h00;
mem[16'hC6FD] = 8'h00;
mem[16'hC6FE] = 8'h00;
mem[16'hC6FF] = 8'h00;
mem[16'hC700] = 8'h00;
mem[16'hC701] = 8'h00;
mem[16'hC702] = 8'h00;
mem[16'hC703] = 8'h00;
mem[16'hC704] = 8'h00;
mem[16'hC705] = 8'h00;
mem[16'hC706] = 8'h00;
mem[16'hC707] = 8'h00;
mem[16'hC708] = 8'h00;
mem[16'hC709] = 8'h00;
mem[16'hC70A] = 8'h00;
mem[16'hC70B] = 8'h00;
mem[16'hC70C] = 8'h00;
mem[16'hC70D] = 8'h00;
mem[16'hC70E] = 8'h00;
mem[16'hC70F] = 8'h00;
mem[16'hC710] = 8'h00;
mem[16'hC711] = 8'h00;
mem[16'hC712] = 8'h00;
mem[16'hC713] = 8'h00;
mem[16'hC714] = 8'h00;
mem[16'hC715] = 8'h00;
mem[16'hC716] = 8'h00;
mem[16'hC717] = 8'h00;
mem[16'hC718] = 8'h00;
mem[16'hC719] = 8'h00;
mem[16'hC71A] = 8'h00;
mem[16'hC71B] = 8'h00;
mem[16'hC71C] = 8'h00;
mem[16'hC71D] = 8'h00;
mem[16'hC71E] = 8'h00;
mem[16'hC71F] = 8'h00;
mem[16'hC720] = 8'h00;
mem[16'hC721] = 8'h00;
mem[16'hC722] = 8'h00;
mem[16'hC723] = 8'h00;
mem[16'hC724] = 8'h00;
mem[16'hC725] = 8'h00;
mem[16'hC726] = 8'h00;
mem[16'hC727] = 8'h00;
mem[16'hC728] = 8'h00;
mem[16'hC729] = 8'h00;
mem[16'hC72A] = 8'h00;
mem[16'hC72B] = 8'h00;
mem[16'hC72C] = 8'h00;
mem[16'hC72D] = 8'h00;
mem[16'hC72E] = 8'h00;
mem[16'hC72F] = 8'h00;
mem[16'hC730] = 8'h00;
mem[16'hC731] = 8'h00;
mem[16'hC732] = 8'h00;
mem[16'hC733] = 8'h00;
mem[16'hC734] = 8'h00;
mem[16'hC735] = 8'h00;
mem[16'hC736] = 8'h00;
mem[16'hC737] = 8'h00;
mem[16'hC738] = 8'h00;
mem[16'hC739] = 8'h00;
mem[16'hC73A] = 8'h00;
mem[16'hC73B] = 8'h00;
mem[16'hC73C] = 8'h00;
mem[16'hC73D] = 8'h00;
mem[16'hC73E] = 8'h00;
mem[16'hC73F] = 8'h00;
mem[16'hC740] = 8'h00;
mem[16'hC741] = 8'h00;
mem[16'hC742] = 8'h00;
mem[16'hC743] = 8'h00;
mem[16'hC744] = 8'h00;
mem[16'hC745] = 8'h00;
mem[16'hC746] = 8'h00;
mem[16'hC747] = 8'h00;
mem[16'hC748] = 8'h00;
mem[16'hC749] = 8'h00;
mem[16'hC74A] = 8'h00;
mem[16'hC74B] = 8'h00;
mem[16'hC74C] = 8'h00;
mem[16'hC74D] = 8'h00;
mem[16'hC74E] = 8'h00;
mem[16'hC74F] = 8'h00;
mem[16'hC750] = 8'h00;
mem[16'hC751] = 8'h00;
mem[16'hC752] = 8'h00;
mem[16'hC753] = 8'h00;
mem[16'hC754] = 8'h00;
mem[16'hC755] = 8'h00;
mem[16'hC756] = 8'h00;
mem[16'hC757] = 8'h00;
mem[16'hC758] = 8'h00;
mem[16'hC759] = 8'h00;
mem[16'hC75A] = 8'h00;
mem[16'hC75B] = 8'h00;
mem[16'hC75C] = 8'h00;
mem[16'hC75D] = 8'h00;
mem[16'hC75E] = 8'h00;
mem[16'hC75F] = 8'h00;
mem[16'hC760] = 8'h00;
mem[16'hC761] = 8'h00;
mem[16'hC762] = 8'h00;
mem[16'hC763] = 8'h00;
mem[16'hC764] = 8'h00;
mem[16'hC765] = 8'h00;
mem[16'hC766] = 8'h00;
mem[16'hC767] = 8'h00;
mem[16'hC768] = 8'h00;
mem[16'hC769] = 8'h00;
mem[16'hC76A] = 8'h00;
mem[16'hC76B] = 8'h00;
mem[16'hC76C] = 8'h00;
mem[16'hC76D] = 8'h00;
mem[16'hC76E] = 8'h00;
mem[16'hC76F] = 8'h00;
mem[16'hC770] = 8'h00;
mem[16'hC771] = 8'h00;
mem[16'hC772] = 8'h00;
mem[16'hC773] = 8'h00;
mem[16'hC774] = 8'h00;
mem[16'hC775] = 8'h00;
mem[16'hC776] = 8'h00;
mem[16'hC777] = 8'h00;
mem[16'hC778] = 8'h00;
mem[16'hC779] = 8'h00;
mem[16'hC77A] = 8'h00;
mem[16'hC77B] = 8'h00;
mem[16'hC77C] = 8'h00;
mem[16'hC77D] = 8'h00;
mem[16'hC77E] = 8'h00;
mem[16'hC77F] = 8'h00;
mem[16'hC780] = 8'h00;
mem[16'hC781] = 8'h00;
mem[16'hC782] = 8'h00;
mem[16'hC783] = 8'h00;
mem[16'hC784] = 8'h00;
mem[16'hC785] = 8'h00;
mem[16'hC786] = 8'h00;
mem[16'hC787] = 8'h00;
mem[16'hC788] = 8'h00;
mem[16'hC789] = 8'h00;
mem[16'hC78A] = 8'h00;
mem[16'hC78B] = 8'h00;
mem[16'hC78C] = 8'h00;
mem[16'hC78D] = 8'h00;
mem[16'hC78E] = 8'h00;
mem[16'hC78F] = 8'h00;
mem[16'hC790] = 8'h00;
mem[16'hC791] = 8'h00;
mem[16'hC792] = 8'h00;
mem[16'hC793] = 8'h00;
mem[16'hC794] = 8'h00;
mem[16'hC795] = 8'h00;
mem[16'hC796] = 8'h00;
mem[16'hC797] = 8'h00;
mem[16'hC798] = 8'h00;
mem[16'hC799] = 8'h00;
mem[16'hC79A] = 8'h00;
mem[16'hC79B] = 8'h00;
mem[16'hC79C] = 8'h00;
mem[16'hC79D] = 8'h00;
mem[16'hC79E] = 8'h00;
mem[16'hC79F] = 8'h00;
mem[16'hC7A0] = 8'h00;
mem[16'hC7A1] = 8'h00;
mem[16'hC7A2] = 8'h00;
mem[16'hC7A3] = 8'h00;
mem[16'hC7A4] = 8'h00;
mem[16'hC7A5] = 8'h00;
mem[16'hC7A6] = 8'h00;
mem[16'hC7A7] = 8'h00;
mem[16'hC7A8] = 8'h00;
mem[16'hC7A9] = 8'h00;
mem[16'hC7AA] = 8'h00;
mem[16'hC7AB] = 8'h00;
mem[16'hC7AC] = 8'h00;
mem[16'hC7AD] = 8'h00;
mem[16'hC7AE] = 8'h00;
mem[16'hC7AF] = 8'h00;
mem[16'hC7B0] = 8'h00;
mem[16'hC7B1] = 8'h00;
mem[16'hC7B2] = 8'h00;
mem[16'hC7B3] = 8'h00;
mem[16'hC7B4] = 8'h00;
mem[16'hC7B5] = 8'h00;
mem[16'hC7B6] = 8'h00;
mem[16'hC7B7] = 8'h00;
mem[16'hC7B8] = 8'h00;
mem[16'hC7B9] = 8'h00;
mem[16'hC7BA] = 8'h00;
mem[16'hC7BB] = 8'h00;
mem[16'hC7BC] = 8'h00;
mem[16'hC7BD] = 8'h00;
mem[16'hC7BE] = 8'h00;
mem[16'hC7BF] = 8'h00;
mem[16'hC7C0] = 8'h00;
mem[16'hC7C1] = 8'h00;
mem[16'hC7C2] = 8'h00;
mem[16'hC7C3] = 8'h00;
mem[16'hC7C4] = 8'h00;
mem[16'hC7C5] = 8'h00;
mem[16'hC7C6] = 8'h00;
mem[16'hC7C7] = 8'h00;
mem[16'hC7C8] = 8'h00;
mem[16'hC7C9] = 8'h00;
mem[16'hC7CA] = 8'h00;
mem[16'hC7CB] = 8'h00;
mem[16'hC7CC] = 8'h00;
mem[16'hC7CD] = 8'h00;
mem[16'hC7CE] = 8'h00;
mem[16'hC7CF] = 8'h00;
mem[16'hC7D0] = 8'h00;
mem[16'hC7D1] = 8'h00;
mem[16'hC7D2] = 8'h00;
mem[16'hC7D3] = 8'h00;
mem[16'hC7D4] = 8'h00;
mem[16'hC7D5] = 8'h00;
mem[16'hC7D6] = 8'h00;
mem[16'hC7D7] = 8'h00;
mem[16'hC7D8] = 8'h00;
mem[16'hC7D9] = 8'h00;
mem[16'hC7DA] = 8'h00;
mem[16'hC7DB] = 8'h00;
mem[16'hC7DC] = 8'h00;
mem[16'hC7DD] = 8'h00;
mem[16'hC7DE] = 8'h00;
mem[16'hC7DF] = 8'h00;
mem[16'hC7E0] = 8'h00;
mem[16'hC7E1] = 8'h00;
mem[16'hC7E2] = 8'h00;
mem[16'hC7E3] = 8'h00;
mem[16'hC7E4] = 8'h00;
mem[16'hC7E5] = 8'h00;
mem[16'hC7E6] = 8'h00;
mem[16'hC7E7] = 8'h00;
mem[16'hC7E8] = 8'h00;
mem[16'hC7E9] = 8'h00;
mem[16'hC7EA] = 8'h00;
mem[16'hC7EB] = 8'h00;
mem[16'hC7EC] = 8'h00;
mem[16'hC7ED] = 8'h00;
mem[16'hC7EE] = 8'h00;
mem[16'hC7EF] = 8'h00;
mem[16'hC7F0] = 8'h00;
mem[16'hC7F1] = 8'h00;
mem[16'hC7F2] = 8'h00;
mem[16'hC7F3] = 8'h00;
mem[16'hC7F4] = 8'h00;
mem[16'hC7F5] = 8'h00;
mem[16'hC7F6] = 8'h00;
mem[16'hC7F7] = 8'h00;
mem[16'hC7F8] = 8'h00;
mem[16'hC7F9] = 8'h00;
mem[16'hC7FA] = 8'h00;
mem[16'hC7FB] = 8'h00;
mem[16'hC7FC] = 8'h00;
mem[16'hC7FD] = 8'h00;
mem[16'hC7FE] = 8'h00;
mem[16'hC7FF] = 8'h00;
mem[16'hC800] = 8'h00;
mem[16'hC801] = 8'h00;
mem[16'hC802] = 8'h00;
mem[16'hC803] = 8'h00;
mem[16'hC804] = 8'h00;
mem[16'hC805] = 8'h00;
mem[16'hC806] = 8'h00;
mem[16'hC807] = 8'h00;
mem[16'hC808] = 8'h00;
mem[16'hC809] = 8'h00;
mem[16'hC80A] = 8'h00;
mem[16'hC80B] = 8'h00;
mem[16'hC80C] = 8'h00;
mem[16'hC80D] = 8'h00;
mem[16'hC80E] = 8'h00;
mem[16'hC80F] = 8'h00;
mem[16'hC810] = 8'h00;
mem[16'hC811] = 8'h00;
mem[16'hC812] = 8'h00;
mem[16'hC813] = 8'h00;
mem[16'hC814] = 8'h00;
mem[16'hC815] = 8'h00;
mem[16'hC816] = 8'h00;
mem[16'hC817] = 8'h00;
mem[16'hC818] = 8'h00;
mem[16'hC819] = 8'h00;
mem[16'hC81A] = 8'h00;
mem[16'hC81B] = 8'h00;
mem[16'hC81C] = 8'h00;
mem[16'hC81D] = 8'h00;
mem[16'hC81E] = 8'h00;
mem[16'hC81F] = 8'h00;
mem[16'hC820] = 8'h00;
mem[16'hC821] = 8'h00;
mem[16'hC822] = 8'h00;
mem[16'hC823] = 8'h00;
mem[16'hC824] = 8'h00;
mem[16'hC825] = 8'h00;
mem[16'hC826] = 8'h00;
mem[16'hC827] = 8'h00;
mem[16'hC828] = 8'h00;
mem[16'hC829] = 8'h00;
mem[16'hC82A] = 8'h00;
mem[16'hC82B] = 8'h00;
mem[16'hC82C] = 8'h00;
mem[16'hC82D] = 8'h00;
mem[16'hC82E] = 8'h00;
mem[16'hC82F] = 8'h00;
mem[16'hC830] = 8'h00;
mem[16'hC831] = 8'h00;
mem[16'hC832] = 8'h00;
mem[16'hC833] = 8'h00;
mem[16'hC834] = 8'h00;
mem[16'hC835] = 8'h00;
mem[16'hC836] = 8'h00;
mem[16'hC837] = 8'h00;
mem[16'hC838] = 8'h00;
mem[16'hC839] = 8'h00;
mem[16'hC83A] = 8'h00;
mem[16'hC83B] = 8'h00;
mem[16'hC83C] = 8'h00;
mem[16'hC83D] = 8'h00;
mem[16'hC83E] = 8'h00;
mem[16'hC83F] = 8'h00;
mem[16'hC840] = 8'h00;
mem[16'hC841] = 8'h00;
mem[16'hC842] = 8'h00;
mem[16'hC843] = 8'h00;
mem[16'hC844] = 8'h00;
mem[16'hC845] = 8'h00;
mem[16'hC846] = 8'h00;
mem[16'hC847] = 8'h00;
mem[16'hC848] = 8'h00;
mem[16'hC849] = 8'h00;
mem[16'hC84A] = 8'h00;
mem[16'hC84B] = 8'h00;
mem[16'hC84C] = 8'h00;
mem[16'hC84D] = 8'h00;
mem[16'hC84E] = 8'h00;
mem[16'hC84F] = 8'h00;
mem[16'hC850] = 8'h00;
mem[16'hC851] = 8'h00;
mem[16'hC852] = 8'h00;
mem[16'hC853] = 8'h00;
mem[16'hC854] = 8'h00;
mem[16'hC855] = 8'h00;
mem[16'hC856] = 8'h00;
mem[16'hC857] = 8'h00;
mem[16'hC858] = 8'h00;
mem[16'hC859] = 8'h00;
mem[16'hC85A] = 8'h00;
mem[16'hC85B] = 8'h00;
mem[16'hC85C] = 8'h00;
mem[16'hC85D] = 8'h00;
mem[16'hC85E] = 8'h00;
mem[16'hC85F] = 8'h00;
mem[16'hC860] = 8'h00;
mem[16'hC861] = 8'h00;
mem[16'hC862] = 8'h00;
mem[16'hC863] = 8'h00;
mem[16'hC864] = 8'h00;
mem[16'hC865] = 8'h00;
mem[16'hC866] = 8'h00;
mem[16'hC867] = 8'h00;
mem[16'hC868] = 8'h00;
mem[16'hC869] = 8'h00;
mem[16'hC86A] = 8'h00;
mem[16'hC86B] = 8'h00;
mem[16'hC86C] = 8'h00;
mem[16'hC86D] = 8'h00;
mem[16'hC86E] = 8'h00;
mem[16'hC86F] = 8'h00;
mem[16'hC870] = 8'h00;
mem[16'hC871] = 8'h00;
mem[16'hC872] = 8'h00;
mem[16'hC873] = 8'h00;
mem[16'hC874] = 8'h00;
mem[16'hC875] = 8'h00;
mem[16'hC876] = 8'h00;
mem[16'hC877] = 8'h00;
mem[16'hC878] = 8'h00;
mem[16'hC879] = 8'h00;
mem[16'hC87A] = 8'h00;
mem[16'hC87B] = 8'h00;
mem[16'hC87C] = 8'h00;
mem[16'hC87D] = 8'h00;
mem[16'hC87E] = 8'h00;
mem[16'hC87F] = 8'h00;
mem[16'hC880] = 8'h00;
mem[16'hC881] = 8'h00;
mem[16'hC882] = 8'h00;
mem[16'hC883] = 8'h00;
mem[16'hC884] = 8'h00;
mem[16'hC885] = 8'h00;
mem[16'hC886] = 8'h00;
mem[16'hC887] = 8'h00;
mem[16'hC888] = 8'h00;
mem[16'hC889] = 8'h00;
mem[16'hC88A] = 8'h00;
mem[16'hC88B] = 8'h00;
mem[16'hC88C] = 8'h00;
mem[16'hC88D] = 8'h00;
mem[16'hC88E] = 8'h00;
mem[16'hC88F] = 8'h00;
mem[16'hC890] = 8'h00;
mem[16'hC891] = 8'h00;
mem[16'hC892] = 8'h00;
mem[16'hC893] = 8'h00;
mem[16'hC894] = 8'h00;
mem[16'hC895] = 8'h00;
mem[16'hC896] = 8'h00;
mem[16'hC897] = 8'h00;
mem[16'hC898] = 8'h00;
mem[16'hC899] = 8'h00;
mem[16'hC89A] = 8'h00;
mem[16'hC89B] = 8'h00;
mem[16'hC89C] = 8'h00;
mem[16'hC89D] = 8'h00;
mem[16'hC89E] = 8'h00;
mem[16'hC89F] = 8'h00;
mem[16'hC8A0] = 8'h00;
mem[16'hC8A1] = 8'h00;
mem[16'hC8A2] = 8'h00;
mem[16'hC8A3] = 8'h00;
mem[16'hC8A4] = 8'h00;
mem[16'hC8A5] = 8'h00;
mem[16'hC8A6] = 8'h00;
mem[16'hC8A7] = 8'h00;
mem[16'hC8A8] = 8'h00;
mem[16'hC8A9] = 8'h00;
mem[16'hC8AA] = 8'h00;
mem[16'hC8AB] = 8'h00;
mem[16'hC8AC] = 8'h00;
mem[16'hC8AD] = 8'h00;
mem[16'hC8AE] = 8'h00;
mem[16'hC8AF] = 8'h00;
mem[16'hC8B0] = 8'h00;
mem[16'hC8B1] = 8'h00;
mem[16'hC8B2] = 8'h00;
mem[16'hC8B3] = 8'h00;
mem[16'hC8B4] = 8'h00;
mem[16'hC8B5] = 8'h00;
mem[16'hC8B6] = 8'h00;
mem[16'hC8B7] = 8'h00;
mem[16'hC8B8] = 8'h00;
mem[16'hC8B9] = 8'h00;
mem[16'hC8BA] = 8'h00;
mem[16'hC8BB] = 8'h00;
mem[16'hC8BC] = 8'h00;
mem[16'hC8BD] = 8'h00;
mem[16'hC8BE] = 8'h00;
mem[16'hC8BF] = 8'h00;
mem[16'hC8C0] = 8'h00;
mem[16'hC8C1] = 8'h00;
mem[16'hC8C2] = 8'h00;
mem[16'hC8C3] = 8'h00;
mem[16'hC8C4] = 8'h00;
mem[16'hC8C5] = 8'h00;
mem[16'hC8C6] = 8'h00;
mem[16'hC8C7] = 8'h00;
mem[16'hC8C8] = 8'h00;
mem[16'hC8C9] = 8'h00;
mem[16'hC8CA] = 8'h00;
mem[16'hC8CB] = 8'h00;
mem[16'hC8CC] = 8'h00;
mem[16'hC8CD] = 8'h00;
mem[16'hC8CE] = 8'h00;
mem[16'hC8CF] = 8'h00;
mem[16'hC8D0] = 8'h00;
mem[16'hC8D1] = 8'h00;
mem[16'hC8D2] = 8'h00;
mem[16'hC8D3] = 8'h00;
mem[16'hC8D4] = 8'h00;
mem[16'hC8D5] = 8'h00;
mem[16'hC8D6] = 8'h00;
mem[16'hC8D7] = 8'h00;
mem[16'hC8D8] = 8'h00;
mem[16'hC8D9] = 8'h00;
mem[16'hC8DA] = 8'h00;
mem[16'hC8DB] = 8'h00;
mem[16'hC8DC] = 8'h00;
mem[16'hC8DD] = 8'h00;
mem[16'hC8DE] = 8'h00;
mem[16'hC8DF] = 8'h00;
mem[16'hC8E0] = 8'h00;
mem[16'hC8E1] = 8'h00;
mem[16'hC8E2] = 8'h00;
mem[16'hC8E3] = 8'h00;
mem[16'hC8E4] = 8'h00;
mem[16'hC8E5] = 8'h00;
mem[16'hC8E6] = 8'h00;
mem[16'hC8E7] = 8'h00;
mem[16'hC8E8] = 8'h00;
mem[16'hC8E9] = 8'h00;
mem[16'hC8EA] = 8'h00;
mem[16'hC8EB] = 8'h00;
mem[16'hC8EC] = 8'h00;
mem[16'hC8ED] = 8'h00;
mem[16'hC8EE] = 8'h00;
mem[16'hC8EF] = 8'h00;
mem[16'hC8F0] = 8'h00;
mem[16'hC8F1] = 8'h00;
mem[16'hC8F2] = 8'h00;
mem[16'hC8F3] = 8'h00;
mem[16'hC8F4] = 8'h00;
mem[16'hC8F5] = 8'h00;
mem[16'hC8F6] = 8'h00;
mem[16'hC8F7] = 8'h00;
mem[16'hC8F8] = 8'h00;
mem[16'hC8F9] = 8'h00;
mem[16'hC8FA] = 8'h00;
mem[16'hC8FB] = 8'h00;
mem[16'hC8FC] = 8'h00;
mem[16'hC8FD] = 8'h00;
mem[16'hC8FE] = 8'h00;
mem[16'hC8FF] = 8'h00;
mem[16'hC900] = 8'h00;
mem[16'hC901] = 8'h00;
mem[16'hC902] = 8'h00;
mem[16'hC903] = 8'h00;
mem[16'hC904] = 8'h00;
mem[16'hC905] = 8'h00;
mem[16'hC906] = 8'h00;
mem[16'hC907] = 8'h00;
mem[16'hC908] = 8'h00;
mem[16'hC909] = 8'h00;
mem[16'hC90A] = 8'h00;
mem[16'hC90B] = 8'h00;
mem[16'hC90C] = 8'h00;
mem[16'hC90D] = 8'h00;
mem[16'hC90E] = 8'h00;
mem[16'hC90F] = 8'h00;
mem[16'hC910] = 8'h00;
mem[16'hC911] = 8'h00;
mem[16'hC912] = 8'h00;
mem[16'hC913] = 8'h00;
mem[16'hC914] = 8'h00;
mem[16'hC915] = 8'h00;
mem[16'hC916] = 8'h00;
mem[16'hC917] = 8'h00;
mem[16'hC918] = 8'h00;
mem[16'hC919] = 8'h00;
mem[16'hC91A] = 8'h00;
mem[16'hC91B] = 8'h00;
mem[16'hC91C] = 8'h00;
mem[16'hC91D] = 8'h00;
mem[16'hC91E] = 8'h00;
mem[16'hC91F] = 8'h00;
mem[16'hC920] = 8'h00;
mem[16'hC921] = 8'h00;
mem[16'hC922] = 8'h00;
mem[16'hC923] = 8'h00;
mem[16'hC924] = 8'h00;
mem[16'hC925] = 8'h00;
mem[16'hC926] = 8'h00;
mem[16'hC927] = 8'h00;
mem[16'hC928] = 8'h00;
mem[16'hC929] = 8'h00;
mem[16'hC92A] = 8'h00;
mem[16'hC92B] = 8'h00;
mem[16'hC92C] = 8'h00;
mem[16'hC92D] = 8'h00;
mem[16'hC92E] = 8'h00;
mem[16'hC92F] = 8'h00;
mem[16'hC930] = 8'h00;
mem[16'hC931] = 8'h00;
mem[16'hC932] = 8'h00;
mem[16'hC933] = 8'h00;
mem[16'hC934] = 8'h00;
mem[16'hC935] = 8'h00;
mem[16'hC936] = 8'h00;
mem[16'hC937] = 8'h00;
mem[16'hC938] = 8'h00;
mem[16'hC939] = 8'h00;
mem[16'hC93A] = 8'h00;
mem[16'hC93B] = 8'h00;
mem[16'hC93C] = 8'h00;
mem[16'hC93D] = 8'h00;
mem[16'hC93E] = 8'h00;
mem[16'hC93F] = 8'h00;
mem[16'hC940] = 8'h00;
mem[16'hC941] = 8'h00;
mem[16'hC942] = 8'h00;
mem[16'hC943] = 8'h00;
mem[16'hC944] = 8'h00;
mem[16'hC945] = 8'h00;
mem[16'hC946] = 8'h00;
mem[16'hC947] = 8'h00;
mem[16'hC948] = 8'h00;
mem[16'hC949] = 8'h00;
mem[16'hC94A] = 8'h00;
mem[16'hC94B] = 8'h00;
mem[16'hC94C] = 8'h00;
mem[16'hC94D] = 8'h00;
mem[16'hC94E] = 8'h00;
mem[16'hC94F] = 8'h00;
mem[16'hC950] = 8'h00;
mem[16'hC951] = 8'h00;
mem[16'hC952] = 8'h00;
mem[16'hC953] = 8'h00;
mem[16'hC954] = 8'h00;
mem[16'hC955] = 8'h00;
mem[16'hC956] = 8'h00;
mem[16'hC957] = 8'h00;
mem[16'hC958] = 8'h00;
mem[16'hC959] = 8'h00;
mem[16'hC95A] = 8'h00;
mem[16'hC95B] = 8'h00;
mem[16'hC95C] = 8'h00;
mem[16'hC95D] = 8'h00;
mem[16'hC95E] = 8'h00;
mem[16'hC95F] = 8'h00;
mem[16'hC960] = 8'h00;
mem[16'hC961] = 8'h00;
mem[16'hC962] = 8'h00;
mem[16'hC963] = 8'h00;
mem[16'hC964] = 8'h00;
mem[16'hC965] = 8'h00;
mem[16'hC966] = 8'h00;
mem[16'hC967] = 8'h00;
mem[16'hC968] = 8'h00;
mem[16'hC969] = 8'h00;
mem[16'hC96A] = 8'h00;
mem[16'hC96B] = 8'h00;
mem[16'hC96C] = 8'h00;
mem[16'hC96D] = 8'h00;
mem[16'hC96E] = 8'h00;
mem[16'hC96F] = 8'h00;
mem[16'hC970] = 8'h00;
mem[16'hC971] = 8'h00;
mem[16'hC972] = 8'h00;
mem[16'hC973] = 8'h00;
mem[16'hC974] = 8'h00;
mem[16'hC975] = 8'h00;
mem[16'hC976] = 8'h00;
mem[16'hC977] = 8'h00;
mem[16'hC978] = 8'h00;
mem[16'hC979] = 8'h00;
mem[16'hC97A] = 8'h00;
mem[16'hC97B] = 8'h00;
mem[16'hC97C] = 8'h00;
mem[16'hC97D] = 8'h00;
mem[16'hC97E] = 8'h00;
mem[16'hC97F] = 8'h00;
mem[16'hC980] = 8'h00;
mem[16'hC981] = 8'h00;
mem[16'hC982] = 8'h00;
mem[16'hC983] = 8'h00;
mem[16'hC984] = 8'h00;
mem[16'hC985] = 8'h00;
mem[16'hC986] = 8'h00;
mem[16'hC987] = 8'h00;
mem[16'hC988] = 8'h00;
mem[16'hC989] = 8'h00;
mem[16'hC98A] = 8'h00;
mem[16'hC98B] = 8'h00;
mem[16'hC98C] = 8'h00;
mem[16'hC98D] = 8'h00;
mem[16'hC98E] = 8'h00;
mem[16'hC98F] = 8'h00;
mem[16'hC990] = 8'h00;
mem[16'hC991] = 8'h00;
mem[16'hC992] = 8'h00;
mem[16'hC993] = 8'h00;
mem[16'hC994] = 8'h00;
mem[16'hC995] = 8'h00;
mem[16'hC996] = 8'h00;
mem[16'hC997] = 8'h00;
mem[16'hC998] = 8'h00;
mem[16'hC999] = 8'h00;
mem[16'hC99A] = 8'h00;
mem[16'hC99B] = 8'h00;
mem[16'hC99C] = 8'h00;
mem[16'hC99D] = 8'h00;
mem[16'hC99E] = 8'h00;
mem[16'hC99F] = 8'h00;
mem[16'hC9A0] = 8'h00;
mem[16'hC9A1] = 8'h00;
mem[16'hC9A2] = 8'h00;
mem[16'hC9A3] = 8'h00;
mem[16'hC9A4] = 8'h00;
mem[16'hC9A5] = 8'h00;
mem[16'hC9A6] = 8'h00;
mem[16'hC9A7] = 8'h00;
mem[16'hC9A8] = 8'h00;
mem[16'hC9A9] = 8'h00;
mem[16'hC9AA] = 8'h00;
mem[16'hC9AB] = 8'h00;
mem[16'hC9AC] = 8'h00;
mem[16'hC9AD] = 8'h00;
mem[16'hC9AE] = 8'h00;
mem[16'hC9AF] = 8'h00;
mem[16'hC9B0] = 8'h00;
mem[16'hC9B1] = 8'h00;
mem[16'hC9B2] = 8'h00;
mem[16'hC9B3] = 8'h00;
mem[16'hC9B4] = 8'h00;
mem[16'hC9B5] = 8'h00;
mem[16'hC9B6] = 8'h00;
mem[16'hC9B7] = 8'h00;
mem[16'hC9B8] = 8'h00;
mem[16'hC9B9] = 8'h00;
mem[16'hC9BA] = 8'h00;
mem[16'hC9BB] = 8'h00;
mem[16'hC9BC] = 8'h00;
mem[16'hC9BD] = 8'h00;
mem[16'hC9BE] = 8'h00;
mem[16'hC9BF] = 8'h00;
mem[16'hC9C0] = 8'h00;
mem[16'hC9C1] = 8'h00;
mem[16'hC9C2] = 8'h00;
mem[16'hC9C3] = 8'h00;
mem[16'hC9C4] = 8'h00;
mem[16'hC9C5] = 8'h00;
mem[16'hC9C6] = 8'h00;
mem[16'hC9C7] = 8'h00;
mem[16'hC9C8] = 8'h00;
mem[16'hC9C9] = 8'h00;
mem[16'hC9CA] = 8'h00;
mem[16'hC9CB] = 8'h00;
mem[16'hC9CC] = 8'h00;
mem[16'hC9CD] = 8'h00;
mem[16'hC9CE] = 8'h00;
mem[16'hC9CF] = 8'h00;
mem[16'hC9D0] = 8'h00;
mem[16'hC9D1] = 8'h00;
mem[16'hC9D2] = 8'h00;
mem[16'hC9D3] = 8'h00;
mem[16'hC9D4] = 8'h00;
mem[16'hC9D5] = 8'h00;
mem[16'hC9D6] = 8'h00;
mem[16'hC9D7] = 8'h00;
mem[16'hC9D8] = 8'h00;
mem[16'hC9D9] = 8'h00;
mem[16'hC9DA] = 8'h00;
mem[16'hC9DB] = 8'h00;
mem[16'hC9DC] = 8'h00;
mem[16'hC9DD] = 8'h00;
mem[16'hC9DE] = 8'h00;
mem[16'hC9DF] = 8'h00;
mem[16'hC9E0] = 8'h00;
mem[16'hC9E1] = 8'h00;
mem[16'hC9E2] = 8'h00;
mem[16'hC9E3] = 8'h00;
mem[16'hC9E4] = 8'h00;
mem[16'hC9E5] = 8'h00;
mem[16'hC9E6] = 8'h00;
mem[16'hC9E7] = 8'h00;
mem[16'hC9E8] = 8'h00;
mem[16'hC9E9] = 8'h00;
mem[16'hC9EA] = 8'h00;
mem[16'hC9EB] = 8'h00;
mem[16'hC9EC] = 8'h00;
mem[16'hC9ED] = 8'h00;
mem[16'hC9EE] = 8'h00;
mem[16'hC9EF] = 8'h00;
mem[16'hC9F0] = 8'h00;
mem[16'hC9F1] = 8'h00;
mem[16'hC9F2] = 8'h00;
mem[16'hC9F3] = 8'h00;
mem[16'hC9F4] = 8'h00;
mem[16'hC9F5] = 8'h00;
mem[16'hC9F6] = 8'h00;
mem[16'hC9F7] = 8'h00;
mem[16'hC9F8] = 8'h00;
mem[16'hC9F9] = 8'h00;
mem[16'hC9FA] = 8'h00;
mem[16'hC9FB] = 8'h00;
mem[16'hC9FC] = 8'h00;
mem[16'hC9FD] = 8'h00;
mem[16'hC9FE] = 8'h00;
mem[16'hC9FF] = 8'h00;
mem[16'hCA00] = 8'h00;
mem[16'hCA01] = 8'h00;
mem[16'hCA02] = 8'h00;
mem[16'hCA03] = 8'h00;
mem[16'hCA04] = 8'h00;
mem[16'hCA05] = 8'h00;
mem[16'hCA06] = 8'h00;
mem[16'hCA07] = 8'h00;
mem[16'hCA08] = 8'h00;
mem[16'hCA09] = 8'h00;
mem[16'hCA0A] = 8'h00;
mem[16'hCA0B] = 8'h00;
mem[16'hCA0C] = 8'h00;
mem[16'hCA0D] = 8'h00;
mem[16'hCA0E] = 8'h00;
mem[16'hCA0F] = 8'h00;
mem[16'hCA10] = 8'h00;
mem[16'hCA11] = 8'h00;
mem[16'hCA12] = 8'h00;
mem[16'hCA13] = 8'h00;
mem[16'hCA14] = 8'h00;
mem[16'hCA15] = 8'h00;
mem[16'hCA16] = 8'h00;
mem[16'hCA17] = 8'h00;
mem[16'hCA18] = 8'h00;
mem[16'hCA19] = 8'h00;
mem[16'hCA1A] = 8'h00;
mem[16'hCA1B] = 8'h00;
mem[16'hCA1C] = 8'h00;
mem[16'hCA1D] = 8'h00;
mem[16'hCA1E] = 8'h00;
mem[16'hCA1F] = 8'h00;
mem[16'hCA20] = 8'h00;
mem[16'hCA21] = 8'h00;
mem[16'hCA22] = 8'h00;
mem[16'hCA23] = 8'h00;
mem[16'hCA24] = 8'h00;
mem[16'hCA25] = 8'h00;
mem[16'hCA26] = 8'h00;
mem[16'hCA27] = 8'h00;
mem[16'hCA28] = 8'h00;
mem[16'hCA29] = 8'h00;
mem[16'hCA2A] = 8'h00;
mem[16'hCA2B] = 8'h00;
mem[16'hCA2C] = 8'h00;
mem[16'hCA2D] = 8'h00;
mem[16'hCA2E] = 8'h00;
mem[16'hCA2F] = 8'h00;
mem[16'hCA30] = 8'h00;
mem[16'hCA31] = 8'h00;
mem[16'hCA32] = 8'h00;
mem[16'hCA33] = 8'h00;
mem[16'hCA34] = 8'h00;
mem[16'hCA35] = 8'h00;
mem[16'hCA36] = 8'h00;
mem[16'hCA37] = 8'h00;
mem[16'hCA38] = 8'h00;
mem[16'hCA39] = 8'h00;
mem[16'hCA3A] = 8'h00;
mem[16'hCA3B] = 8'h00;
mem[16'hCA3C] = 8'h00;
mem[16'hCA3D] = 8'h00;
mem[16'hCA3E] = 8'h00;
mem[16'hCA3F] = 8'h00;
mem[16'hCA40] = 8'h00;
mem[16'hCA41] = 8'h00;
mem[16'hCA42] = 8'h00;
mem[16'hCA43] = 8'h00;
mem[16'hCA44] = 8'h00;
mem[16'hCA45] = 8'h00;
mem[16'hCA46] = 8'h00;
mem[16'hCA47] = 8'h00;
mem[16'hCA48] = 8'h00;
mem[16'hCA49] = 8'h00;
mem[16'hCA4A] = 8'h00;
mem[16'hCA4B] = 8'h00;
mem[16'hCA4C] = 8'h00;
mem[16'hCA4D] = 8'h00;
mem[16'hCA4E] = 8'h00;
mem[16'hCA4F] = 8'h00;
mem[16'hCA50] = 8'h00;
mem[16'hCA51] = 8'h00;
mem[16'hCA52] = 8'h00;
mem[16'hCA53] = 8'h00;
mem[16'hCA54] = 8'h00;
mem[16'hCA55] = 8'h00;
mem[16'hCA56] = 8'h00;
mem[16'hCA57] = 8'h00;
mem[16'hCA58] = 8'h00;
mem[16'hCA59] = 8'h00;
mem[16'hCA5A] = 8'h00;
mem[16'hCA5B] = 8'h00;
mem[16'hCA5C] = 8'h00;
mem[16'hCA5D] = 8'h00;
mem[16'hCA5E] = 8'h00;
mem[16'hCA5F] = 8'h00;
mem[16'hCA60] = 8'h00;
mem[16'hCA61] = 8'h00;
mem[16'hCA62] = 8'h00;
mem[16'hCA63] = 8'h00;
mem[16'hCA64] = 8'h00;
mem[16'hCA65] = 8'h00;
mem[16'hCA66] = 8'h00;
mem[16'hCA67] = 8'h00;
mem[16'hCA68] = 8'h00;
mem[16'hCA69] = 8'h00;
mem[16'hCA6A] = 8'h00;
mem[16'hCA6B] = 8'h00;
mem[16'hCA6C] = 8'h00;
mem[16'hCA6D] = 8'h00;
mem[16'hCA6E] = 8'h00;
mem[16'hCA6F] = 8'h00;
mem[16'hCA70] = 8'h00;
mem[16'hCA71] = 8'h00;
mem[16'hCA72] = 8'h00;
mem[16'hCA73] = 8'h00;
mem[16'hCA74] = 8'h00;
mem[16'hCA75] = 8'h00;
mem[16'hCA76] = 8'h00;
mem[16'hCA77] = 8'h00;
mem[16'hCA78] = 8'h00;
mem[16'hCA79] = 8'h00;
mem[16'hCA7A] = 8'h00;
mem[16'hCA7B] = 8'h00;
mem[16'hCA7C] = 8'h00;
mem[16'hCA7D] = 8'h00;
mem[16'hCA7E] = 8'h00;
mem[16'hCA7F] = 8'h00;
mem[16'hCA80] = 8'h00;
mem[16'hCA81] = 8'h00;
mem[16'hCA82] = 8'h00;
mem[16'hCA83] = 8'h00;
mem[16'hCA84] = 8'h00;
mem[16'hCA85] = 8'h00;
mem[16'hCA86] = 8'h00;
mem[16'hCA87] = 8'h00;
mem[16'hCA88] = 8'h00;
mem[16'hCA89] = 8'h00;
mem[16'hCA8A] = 8'h00;
mem[16'hCA8B] = 8'h00;
mem[16'hCA8C] = 8'h00;
mem[16'hCA8D] = 8'h00;
mem[16'hCA8E] = 8'h00;
mem[16'hCA8F] = 8'h00;
mem[16'hCA90] = 8'h00;
mem[16'hCA91] = 8'h00;
mem[16'hCA92] = 8'h00;
mem[16'hCA93] = 8'h00;
mem[16'hCA94] = 8'h00;
mem[16'hCA95] = 8'h00;
mem[16'hCA96] = 8'h00;
mem[16'hCA97] = 8'h00;
mem[16'hCA98] = 8'h00;
mem[16'hCA99] = 8'h00;
mem[16'hCA9A] = 8'h00;
mem[16'hCA9B] = 8'h00;
mem[16'hCA9C] = 8'h00;
mem[16'hCA9D] = 8'h00;
mem[16'hCA9E] = 8'h00;
mem[16'hCA9F] = 8'h00;
mem[16'hCAA0] = 8'h00;
mem[16'hCAA1] = 8'h00;
mem[16'hCAA2] = 8'h00;
mem[16'hCAA3] = 8'h00;
mem[16'hCAA4] = 8'h00;
mem[16'hCAA5] = 8'h00;
mem[16'hCAA6] = 8'h00;
mem[16'hCAA7] = 8'h00;
mem[16'hCAA8] = 8'h00;
mem[16'hCAA9] = 8'h00;
mem[16'hCAAA] = 8'h00;
mem[16'hCAAB] = 8'h00;
mem[16'hCAAC] = 8'h00;
mem[16'hCAAD] = 8'h00;
mem[16'hCAAE] = 8'h00;
mem[16'hCAAF] = 8'h00;
mem[16'hCAB0] = 8'h00;
mem[16'hCAB1] = 8'h00;
mem[16'hCAB2] = 8'h00;
mem[16'hCAB3] = 8'h00;
mem[16'hCAB4] = 8'h00;
mem[16'hCAB5] = 8'h00;
mem[16'hCAB6] = 8'h00;
mem[16'hCAB7] = 8'h00;
mem[16'hCAB8] = 8'h00;
mem[16'hCAB9] = 8'h00;
mem[16'hCABA] = 8'h00;
mem[16'hCABB] = 8'h00;
mem[16'hCABC] = 8'h00;
mem[16'hCABD] = 8'h00;
mem[16'hCABE] = 8'h00;
mem[16'hCABF] = 8'h00;
mem[16'hCAC0] = 8'h00;
mem[16'hCAC1] = 8'h00;
mem[16'hCAC2] = 8'h00;
mem[16'hCAC3] = 8'h00;
mem[16'hCAC4] = 8'h00;
mem[16'hCAC5] = 8'h00;
mem[16'hCAC6] = 8'h00;
mem[16'hCAC7] = 8'h00;
mem[16'hCAC8] = 8'h00;
mem[16'hCAC9] = 8'h00;
mem[16'hCACA] = 8'h00;
mem[16'hCACB] = 8'h00;
mem[16'hCACC] = 8'h00;
mem[16'hCACD] = 8'h00;
mem[16'hCACE] = 8'h00;
mem[16'hCACF] = 8'h00;
mem[16'hCAD0] = 8'h00;
mem[16'hCAD1] = 8'h00;
mem[16'hCAD2] = 8'h00;
mem[16'hCAD3] = 8'h00;
mem[16'hCAD4] = 8'h00;
mem[16'hCAD5] = 8'h00;
mem[16'hCAD6] = 8'h00;
mem[16'hCAD7] = 8'h00;
mem[16'hCAD8] = 8'h00;
mem[16'hCAD9] = 8'h00;
mem[16'hCADA] = 8'h00;
mem[16'hCADB] = 8'h00;
mem[16'hCADC] = 8'h00;
mem[16'hCADD] = 8'h00;
mem[16'hCADE] = 8'h00;
mem[16'hCADF] = 8'h00;
mem[16'hCAE0] = 8'h00;
mem[16'hCAE1] = 8'h00;
mem[16'hCAE2] = 8'h00;
mem[16'hCAE3] = 8'h00;
mem[16'hCAE4] = 8'h00;
mem[16'hCAE5] = 8'h00;
mem[16'hCAE6] = 8'h00;
mem[16'hCAE7] = 8'h00;
mem[16'hCAE8] = 8'h00;
mem[16'hCAE9] = 8'h00;
mem[16'hCAEA] = 8'h00;
mem[16'hCAEB] = 8'h00;
mem[16'hCAEC] = 8'h00;
mem[16'hCAED] = 8'h00;
mem[16'hCAEE] = 8'h00;
mem[16'hCAEF] = 8'h00;
mem[16'hCAF0] = 8'h00;
mem[16'hCAF1] = 8'h00;
mem[16'hCAF2] = 8'h00;
mem[16'hCAF3] = 8'h00;
mem[16'hCAF4] = 8'h00;
mem[16'hCAF5] = 8'h00;
mem[16'hCAF6] = 8'h00;
mem[16'hCAF7] = 8'h00;
mem[16'hCAF8] = 8'h00;
mem[16'hCAF9] = 8'h00;
mem[16'hCAFA] = 8'h00;
mem[16'hCAFB] = 8'h00;
mem[16'hCAFC] = 8'h00;
mem[16'hCAFD] = 8'h00;
mem[16'hCAFE] = 8'h00;
mem[16'hCAFF] = 8'h00;
mem[16'hCB00] = 8'h00;
mem[16'hCB01] = 8'h00;
mem[16'hCB02] = 8'h00;
mem[16'hCB03] = 8'h00;
mem[16'hCB04] = 8'h00;
mem[16'hCB05] = 8'h00;
mem[16'hCB06] = 8'h00;
mem[16'hCB07] = 8'h00;
mem[16'hCB08] = 8'h00;
mem[16'hCB09] = 8'h00;
mem[16'hCB0A] = 8'h00;
mem[16'hCB0B] = 8'h00;
mem[16'hCB0C] = 8'h00;
mem[16'hCB0D] = 8'h00;
mem[16'hCB0E] = 8'h00;
mem[16'hCB0F] = 8'h00;
mem[16'hCB10] = 8'h00;
mem[16'hCB11] = 8'h00;
mem[16'hCB12] = 8'h00;
mem[16'hCB13] = 8'h00;
mem[16'hCB14] = 8'h00;
mem[16'hCB15] = 8'h00;
mem[16'hCB16] = 8'h00;
mem[16'hCB17] = 8'h00;
mem[16'hCB18] = 8'h00;
mem[16'hCB19] = 8'h00;
mem[16'hCB1A] = 8'h00;
mem[16'hCB1B] = 8'h00;
mem[16'hCB1C] = 8'h00;
mem[16'hCB1D] = 8'h00;
mem[16'hCB1E] = 8'h00;
mem[16'hCB1F] = 8'h00;
mem[16'hCB20] = 8'h00;
mem[16'hCB21] = 8'h00;
mem[16'hCB22] = 8'h00;
mem[16'hCB23] = 8'h00;
mem[16'hCB24] = 8'h00;
mem[16'hCB25] = 8'h00;
mem[16'hCB26] = 8'h00;
mem[16'hCB27] = 8'h00;
mem[16'hCB28] = 8'h00;
mem[16'hCB29] = 8'h00;
mem[16'hCB2A] = 8'h00;
mem[16'hCB2B] = 8'h00;
mem[16'hCB2C] = 8'h00;
mem[16'hCB2D] = 8'h00;
mem[16'hCB2E] = 8'h00;
mem[16'hCB2F] = 8'h00;
mem[16'hCB30] = 8'h00;
mem[16'hCB31] = 8'h00;
mem[16'hCB32] = 8'h00;
mem[16'hCB33] = 8'h00;
mem[16'hCB34] = 8'h00;
mem[16'hCB35] = 8'h00;
mem[16'hCB36] = 8'h00;
mem[16'hCB37] = 8'h00;
mem[16'hCB38] = 8'h00;
mem[16'hCB39] = 8'h00;
mem[16'hCB3A] = 8'h00;
mem[16'hCB3B] = 8'h00;
mem[16'hCB3C] = 8'h00;
mem[16'hCB3D] = 8'h00;
mem[16'hCB3E] = 8'h00;
mem[16'hCB3F] = 8'h00;
mem[16'hCB40] = 8'h00;
mem[16'hCB41] = 8'h00;
mem[16'hCB42] = 8'h00;
mem[16'hCB43] = 8'h00;
mem[16'hCB44] = 8'h00;
mem[16'hCB45] = 8'h00;
mem[16'hCB46] = 8'h00;
mem[16'hCB47] = 8'h00;
mem[16'hCB48] = 8'h00;
mem[16'hCB49] = 8'h00;
mem[16'hCB4A] = 8'h00;
mem[16'hCB4B] = 8'h00;
mem[16'hCB4C] = 8'h00;
mem[16'hCB4D] = 8'h00;
mem[16'hCB4E] = 8'h00;
mem[16'hCB4F] = 8'h00;
mem[16'hCB50] = 8'h00;
mem[16'hCB51] = 8'h00;
mem[16'hCB52] = 8'h00;
mem[16'hCB53] = 8'h00;
mem[16'hCB54] = 8'h00;
mem[16'hCB55] = 8'h00;
mem[16'hCB56] = 8'h00;
mem[16'hCB57] = 8'h00;
mem[16'hCB58] = 8'h00;
mem[16'hCB59] = 8'h00;
mem[16'hCB5A] = 8'h00;
mem[16'hCB5B] = 8'h00;
mem[16'hCB5C] = 8'h00;
mem[16'hCB5D] = 8'h00;
mem[16'hCB5E] = 8'h00;
mem[16'hCB5F] = 8'h00;
mem[16'hCB60] = 8'h00;
mem[16'hCB61] = 8'h00;
mem[16'hCB62] = 8'h00;
mem[16'hCB63] = 8'h00;
mem[16'hCB64] = 8'h00;
mem[16'hCB65] = 8'h00;
mem[16'hCB66] = 8'h00;
mem[16'hCB67] = 8'h00;
mem[16'hCB68] = 8'h00;
mem[16'hCB69] = 8'h00;
mem[16'hCB6A] = 8'h00;
mem[16'hCB6B] = 8'h00;
mem[16'hCB6C] = 8'h00;
mem[16'hCB6D] = 8'h00;
mem[16'hCB6E] = 8'h00;
mem[16'hCB6F] = 8'h00;
mem[16'hCB70] = 8'h00;
mem[16'hCB71] = 8'h00;
mem[16'hCB72] = 8'h00;
mem[16'hCB73] = 8'h00;
mem[16'hCB74] = 8'h00;
mem[16'hCB75] = 8'h00;
mem[16'hCB76] = 8'h00;
mem[16'hCB77] = 8'h00;
mem[16'hCB78] = 8'h00;
mem[16'hCB79] = 8'h00;
mem[16'hCB7A] = 8'h00;
mem[16'hCB7B] = 8'h00;
mem[16'hCB7C] = 8'h00;
mem[16'hCB7D] = 8'h00;
mem[16'hCB7E] = 8'h00;
mem[16'hCB7F] = 8'h00;
mem[16'hCB80] = 8'h00;
mem[16'hCB81] = 8'h00;
mem[16'hCB82] = 8'h00;
mem[16'hCB83] = 8'h00;
mem[16'hCB84] = 8'h00;
mem[16'hCB85] = 8'h00;
mem[16'hCB86] = 8'h00;
mem[16'hCB87] = 8'h00;
mem[16'hCB88] = 8'h00;
mem[16'hCB89] = 8'h00;
mem[16'hCB8A] = 8'h00;
mem[16'hCB8B] = 8'h00;
mem[16'hCB8C] = 8'h00;
mem[16'hCB8D] = 8'h00;
mem[16'hCB8E] = 8'h00;
mem[16'hCB8F] = 8'h00;
mem[16'hCB90] = 8'h00;
mem[16'hCB91] = 8'h00;
mem[16'hCB92] = 8'h00;
mem[16'hCB93] = 8'h00;
mem[16'hCB94] = 8'h00;
mem[16'hCB95] = 8'h00;
mem[16'hCB96] = 8'h00;
mem[16'hCB97] = 8'h00;
mem[16'hCB98] = 8'h00;
mem[16'hCB99] = 8'h00;
mem[16'hCB9A] = 8'h00;
mem[16'hCB9B] = 8'h00;
mem[16'hCB9C] = 8'h00;
mem[16'hCB9D] = 8'h00;
mem[16'hCB9E] = 8'h00;
mem[16'hCB9F] = 8'h00;
mem[16'hCBA0] = 8'h00;
mem[16'hCBA1] = 8'h00;
mem[16'hCBA2] = 8'h00;
mem[16'hCBA3] = 8'h00;
mem[16'hCBA4] = 8'h00;
mem[16'hCBA5] = 8'h00;
mem[16'hCBA6] = 8'h00;
mem[16'hCBA7] = 8'h00;
mem[16'hCBA8] = 8'h00;
mem[16'hCBA9] = 8'h00;
mem[16'hCBAA] = 8'h00;
mem[16'hCBAB] = 8'h00;
mem[16'hCBAC] = 8'h00;
mem[16'hCBAD] = 8'h00;
mem[16'hCBAE] = 8'h00;
mem[16'hCBAF] = 8'h00;
mem[16'hCBB0] = 8'h00;
mem[16'hCBB1] = 8'h00;
mem[16'hCBB2] = 8'h00;
mem[16'hCBB3] = 8'h00;
mem[16'hCBB4] = 8'h00;
mem[16'hCBB5] = 8'h00;
mem[16'hCBB6] = 8'h00;
mem[16'hCBB7] = 8'h00;
mem[16'hCBB8] = 8'h00;
mem[16'hCBB9] = 8'h00;
mem[16'hCBBA] = 8'h00;
mem[16'hCBBB] = 8'h00;
mem[16'hCBBC] = 8'h00;
mem[16'hCBBD] = 8'h00;
mem[16'hCBBE] = 8'h00;
mem[16'hCBBF] = 8'h00;
mem[16'hCBC0] = 8'h00;
mem[16'hCBC1] = 8'h00;
mem[16'hCBC2] = 8'h00;
mem[16'hCBC3] = 8'h00;
mem[16'hCBC4] = 8'h00;
mem[16'hCBC5] = 8'h00;
mem[16'hCBC6] = 8'h00;
mem[16'hCBC7] = 8'h00;
mem[16'hCBC8] = 8'h00;
mem[16'hCBC9] = 8'h00;
mem[16'hCBCA] = 8'h00;
mem[16'hCBCB] = 8'h00;
mem[16'hCBCC] = 8'h00;
mem[16'hCBCD] = 8'h00;
mem[16'hCBCE] = 8'h00;
mem[16'hCBCF] = 8'h00;
mem[16'hCBD0] = 8'h00;
mem[16'hCBD1] = 8'h00;
mem[16'hCBD2] = 8'h00;
mem[16'hCBD3] = 8'h00;
mem[16'hCBD4] = 8'h00;
mem[16'hCBD5] = 8'h00;
mem[16'hCBD6] = 8'h00;
mem[16'hCBD7] = 8'h00;
mem[16'hCBD8] = 8'h00;
mem[16'hCBD9] = 8'h00;
mem[16'hCBDA] = 8'h00;
mem[16'hCBDB] = 8'h00;
mem[16'hCBDC] = 8'h00;
mem[16'hCBDD] = 8'h00;
mem[16'hCBDE] = 8'h00;
mem[16'hCBDF] = 8'h00;
mem[16'hCBE0] = 8'h00;
mem[16'hCBE1] = 8'h00;
mem[16'hCBE2] = 8'h00;
mem[16'hCBE3] = 8'h00;
mem[16'hCBE4] = 8'h00;
mem[16'hCBE5] = 8'h00;
mem[16'hCBE6] = 8'h00;
mem[16'hCBE7] = 8'h00;
mem[16'hCBE8] = 8'h00;
mem[16'hCBE9] = 8'h00;
mem[16'hCBEA] = 8'h00;
mem[16'hCBEB] = 8'h00;
mem[16'hCBEC] = 8'h00;
mem[16'hCBED] = 8'h00;
mem[16'hCBEE] = 8'h00;
mem[16'hCBEF] = 8'h00;
mem[16'hCBF0] = 8'h00;
mem[16'hCBF1] = 8'h00;
mem[16'hCBF2] = 8'h00;
mem[16'hCBF3] = 8'h00;
mem[16'hCBF4] = 8'h00;
mem[16'hCBF5] = 8'h00;
mem[16'hCBF6] = 8'h00;
mem[16'hCBF7] = 8'h00;
mem[16'hCBF8] = 8'h00;
mem[16'hCBF9] = 8'h00;
mem[16'hCBFA] = 8'h00;
mem[16'hCBFB] = 8'h00;
mem[16'hCBFC] = 8'h00;
mem[16'hCBFD] = 8'h00;
mem[16'hCBFE] = 8'h00;
mem[16'hCBFF] = 8'h00;
mem[16'hCC00] = 8'h00;
mem[16'hCC01] = 8'h00;
mem[16'hCC02] = 8'h00;
mem[16'hCC03] = 8'h00;
mem[16'hCC04] = 8'h00;
mem[16'hCC05] = 8'h00;
mem[16'hCC06] = 8'h00;
mem[16'hCC07] = 8'h00;
mem[16'hCC08] = 8'h00;
mem[16'hCC09] = 8'h00;
mem[16'hCC0A] = 8'h00;
mem[16'hCC0B] = 8'h00;
mem[16'hCC0C] = 8'h00;
mem[16'hCC0D] = 8'h00;
mem[16'hCC0E] = 8'h00;
mem[16'hCC0F] = 8'h00;
mem[16'hCC10] = 8'h00;
mem[16'hCC11] = 8'h00;
mem[16'hCC12] = 8'h00;
mem[16'hCC13] = 8'h00;
mem[16'hCC14] = 8'h00;
mem[16'hCC15] = 8'h00;
mem[16'hCC16] = 8'h00;
mem[16'hCC17] = 8'h00;
mem[16'hCC18] = 8'h00;
mem[16'hCC19] = 8'h00;
mem[16'hCC1A] = 8'h00;
mem[16'hCC1B] = 8'h00;
mem[16'hCC1C] = 8'h00;
mem[16'hCC1D] = 8'h00;
mem[16'hCC1E] = 8'h00;
mem[16'hCC1F] = 8'h00;
mem[16'hCC20] = 8'h00;
mem[16'hCC21] = 8'h00;
mem[16'hCC22] = 8'h00;
mem[16'hCC23] = 8'h00;
mem[16'hCC24] = 8'h00;
mem[16'hCC25] = 8'h00;
mem[16'hCC26] = 8'h00;
mem[16'hCC27] = 8'h00;
mem[16'hCC28] = 8'h00;
mem[16'hCC29] = 8'h00;
mem[16'hCC2A] = 8'h00;
mem[16'hCC2B] = 8'h00;
mem[16'hCC2C] = 8'h00;
mem[16'hCC2D] = 8'h00;
mem[16'hCC2E] = 8'h00;
mem[16'hCC2F] = 8'h00;
mem[16'hCC30] = 8'h00;
mem[16'hCC31] = 8'h00;
mem[16'hCC32] = 8'h00;
mem[16'hCC33] = 8'h00;
mem[16'hCC34] = 8'h00;
mem[16'hCC35] = 8'h00;
mem[16'hCC36] = 8'h00;
mem[16'hCC37] = 8'h00;
mem[16'hCC38] = 8'h00;
mem[16'hCC39] = 8'h00;
mem[16'hCC3A] = 8'h00;
mem[16'hCC3B] = 8'h00;
mem[16'hCC3C] = 8'h00;
mem[16'hCC3D] = 8'h00;
mem[16'hCC3E] = 8'h00;
mem[16'hCC3F] = 8'h00;
mem[16'hCC40] = 8'h00;
mem[16'hCC41] = 8'h00;
mem[16'hCC42] = 8'h00;
mem[16'hCC43] = 8'h00;
mem[16'hCC44] = 8'h00;
mem[16'hCC45] = 8'h00;
mem[16'hCC46] = 8'h00;
mem[16'hCC47] = 8'h00;
mem[16'hCC48] = 8'h00;
mem[16'hCC49] = 8'h00;
mem[16'hCC4A] = 8'h00;
mem[16'hCC4B] = 8'h00;
mem[16'hCC4C] = 8'h00;
mem[16'hCC4D] = 8'h00;
mem[16'hCC4E] = 8'h00;
mem[16'hCC4F] = 8'h00;
mem[16'hCC50] = 8'h00;
mem[16'hCC51] = 8'h00;
mem[16'hCC52] = 8'h00;
mem[16'hCC53] = 8'h00;
mem[16'hCC54] = 8'h00;
mem[16'hCC55] = 8'h00;
mem[16'hCC56] = 8'h00;
mem[16'hCC57] = 8'h00;
mem[16'hCC58] = 8'h00;
mem[16'hCC59] = 8'h00;
mem[16'hCC5A] = 8'h00;
mem[16'hCC5B] = 8'h00;
mem[16'hCC5C] = 8'h00;
mem[16'hCC5D] = 8'h00;
mem[16'hCC5E] = 8'h00;
mem[16'hCC5F] = 8'h00;
mem[16'hCC60] = 8'h00;
mem[16'hCC61] = 8'h00;
mem[16'hCC62] = 8'h00;
mem[16'hCC63] = 8'h00;
mem[16'hCC64] = 8'h00;
mem[16'hCC65] = 8'h00;
mem[16'hCC66] = 8'h00;
mem[16'hCC67] = 8'h00;
mem[16'hCC68] = 8'h00;
mem[16'hCC69] = 8'h00;
mem[16'hCC6A] = 8'h00;
mem[16'hCC6B] = 8'h00;
mem[16'hCC6C] = 8'h00;
mem[16'hCC6D] = 8'h00;
mem[16'hCC6E] = 8'h00;
mem[16'hCC6F] = 8'h00;
mem[16'hCC70] = 8'h00;
mem[16'hCC71] = 8'h00;
mem[16'hCC72] = 8'h00;
mem[16'hCC73] = 8'h00;
mem[16'hCC74] = 8'h00;
mem[16'hCC75] = 8'h00;
mem[16'hCC76] = 8'h00;
mem[16'hCC77] = 8'h00;
mem[16'hCC78] = 8'h00;
mem[16'hCC79] = 8'h00;
mem[16'hCC7A] = 8'h00;
mem[16'hCC7B] = 8'h00;
mem[16'hCC7C] = 8'h00;
mem[16'hCC7D] = 8'h00;
mem[16'hCC7E] = 8'h00;
mem[16'hCC7F] = 8'h00;
mem[16'hCC80] = 8'h00;
mem[16'hCC81] = 8'h00;
mem[16'hCC82] = 8'h00;
mem[16'hCC83] = 8'h00;
mem[16'hCC84] = 8'h00;
mem[16'hCC85] = 8'h00;
mem[16'hCC86] = 8'h00;
mem[16'hCC87] = 8'h00;
mem[16'hCC88] = 8'h00;
mem[16'hCC89] = 8'h00;
mem[16'hCC8A] = 8'h00;
mem[16'hCC8B] = 8'h00;
mem[16'hCC8C] = 8'h00;
mem[16'hCC8D] = 8'h00;
mem[16'hCC8E] = 8'h00;
mem[16'hCC8F] = 8'h00;
mem[16'hCC90] = 8'h00;
mem[16'hCC91] = 8'h00;
mem[16'hCC92] = 8'h00;
mem[16'hCC93] = 8'h00;
mem[16'hCC94] = 8'h00;
mem[16'hCC95] = 8'h00;
mem[16'hCC96] = 8'h00;
mem[16'hCC97] = 8'h00;
mem[16'hCC98] = 8'h00;
mem[16'hCC99] = 8'h00;
mem[16'hCC9A] = 8'h00;
mem[16'hCC9B] = 8'h00;
mem[16'hCC9C] = 8'h00;
mem[16'hCC9D] = 8'h00;
mem[16'hCC9E] = 8'h00;
mem[16'hCC9F] = 8'h00;
mem[16'hCCA0] = 8'h00;
mem[16'hCCA1] = 8'h00;
mem[16'hCCA2] = 8'h00;
mem[16'hCCA3] = 8'h00;
mem[16'hCCA4] = 8'h00;
mem[16'hCCA5] = 8'h00;
mem[16'hCCA6] = 8'h00;
mem[16'hCCA7] = 8'h00;
mem[16'hCCA8] = 8'h00;
mem[16'hCCA9] = 8'h00;
mem[16'hCCAA] = 8'h00;
mem[16'hCCAB] = 8'h00;
mem[16'hCCAC] = 8'h00;
mem[16'hCCAD] = 8'h00;
mem[16'hCCAE] = 8'h00;
mem[16'hCCAF] = 8'h00;
mem[16'hCCB0] = 8'h00;
mem[16'hCCB1] = 8'h00;
mem[16'hCCB2] = 8'h00;
mem[16'hCCB3] = 8'h00;
mem[16'hCCB4] = 8'h00;
mem[16'hCCB5] = 8'h00;
mem[16'hCCB6] = 8'h00;
mem[16'hCCB7] = 8'h00;
mem[16'hCCB8] = 8'h00;
mem[16'hCCB9] = 8'h00;
mem[16'hCCBA] = 8'h00;
mem[16'hCCBB] = 8'h00;
mem[16'hCCBC] = 8'h00;
mem[16'hCCBD] = 8'h00;
mem[16'hCCBE] = 8'h00;
mem[16'hCCBF] = 8'h00;
mem[16'hCCC0] = 8'h00;
mem[16'hCCC1] = 8'h00;
mem[16'hCCC2] = 8'h00;
mem[16'hCCC3] = 8'h00;
mem[16'hCCC4] = 8'h00;
mem[16'hCCC5] = 8'h00;
mem[16'hCCC6] = 8'h00;
mem[16'hCCC7] = 8'h00;
mem[16'hCCC8] = 8'h00;
mem[16'hCCC9] = 8'h00;
mem[16'hCCCA] = 8'h00;
mem[16'hCCCB] = 8'h00;
mem[16'hCCCC] = 8'h00;
mem[16'hCCCD] = 8'h00;
mem[16'hCCCE] = 8'h00;
mem[16'hCCCF] = 8'h00;
mem[16'hCCD0] = 8'h00;
mem[16'hCCD1] = 8'h00;
mem[16'hCCD2] = 8'h00;
mem[16'hCCD3] = 8'h00;
mem[16'hCCD4] = 8'h00;
mem[16'hCCD5] = 8'h00;
mem[16'hCCD6] = 8'h00;
mem[16'hCCD7] = 8'h00;
mem[16'hCCD8] = 8'h00;
mem[16'hCCD9] = 8'h00;
mem[16'hCCDA] = 8'h00;
mem[16'hCCDB] = 8'h00;
mem[16'hCCDC] = 8'h00;
mem[16'hCCDD] = 8'h00;
mem[16'hCCDE] = 8'h00;
mem[16'hCCDF] = 8'h00;
mem[16'hCCE0] = 8'h00;
mem[16'hCCE1] = 8'h00;
mem[16'hCCE2] = 8'h00;
mem[16'hCCE3] = 8'h00;
mem[16'hCCE4] = 8'h00;
mem[16'hCCE5] = 8'h00;
mem[16'hCCE6] = 8'h00;
mem[16'hCCE7] = 8'h00;
mem[16'hCCE8] = 8'h00;
mem[16'hCCE9] = 8'h00;
mem[16'hCCEA] = 8'h00;
mem[16'hCCEB] = 8'h00;
mem[16'hCCEC] = 8'h00;
mem[16'hCCED] = 8'h00;
mem[16'hCCEE] = 8'h00;
mem[16'hCCEF] = 8'h00;
mem[16'hCCF0] = 8'h00;
mem[16'hCCF1] = 8'h00;
mem[16'hCCF2] = 8'h00;
mem[16'hCCF3] = 8'h00;
mem[16'hCCF4] = 8'h00;
mem[16'hCCF5] = 8'h00;
mem[16'hCCF6] = 8'h00;
mem[16'hCCF7] = 8'h00;
mem[16'hCCF8] = 8'h00;
mem[16'hCCF9] = 8'h00;
mem[16'hCCFA] = 8'h00;
mem[16'hCCFB] = 8'h00;
mem[16'hCCFC] = 8'h00;
mem[16'hCCFD] = 8'h00;
mem[16'hCCFE] = 8'h00;
mem[16'hCCFF] = 8'h00;
mem[16'hCD00] = 8'h00;
mem[16'hCD01] = 8'h00;
mem[16'hCD02] = 8'h00;
mem[16'hCD03] = 8'h00;
mem[16'hCD04] = 8'h00;
mem[16'hCD05] = 8'h00;
mem[16'hCD06] = 8'h00;
mem[16'hCD07] = 8'h00;
mem[16'hCD08] = 8'h00;
mem[16'hCD09] = 8'h00;
mem[16'hCD0A] = 8'h00;
mem[16'hCD0B] = 8'h00;
mem[16'hCD0C] = 8'h00;
mem[16'hCD0D] = 8'h00;
mem[16'hCD0E] = 8'h00;
mem[16'hCD0F] = 8'h00;
mem[16'hCD10] = 8'h00;
mem[16'hCD11] = 8'h00;
mem[16'hCD12] = 8'h00;
mem[16'hCD13] = 8'h00;
mem[16'hCD14] = 8'h00;
mem[16'hCD15] = 8'h00;
mem[16'hCD16] = 8'h00;
mem[16'hCD17] = 8'h00;
mem[16'hCD18] = 8'h00;
mem[16'hCD19] = 8'h00;
mem[16'hCD1A] = 8'h00;
mem[16'hCD1B] = 8'h00;
mem[16'hCD1C] = 8'h00;
mem[16'hCD1D] = 8'h00;
mem[16'hCD1E] = 8'h00;
mem[16'hCD1F] = 8'h00;
mem[16'hCD20] = 8'h00;
mem[16'hCD21] = 8'h00;
mem[16'hCD22] = 8'h00;
mem[16'hCD23] = 8'h00;
mem[16'hCD24] = 8'h00;
mem[16'hCD25] = 8'h00;
mem[16'hCD26] = 8'h00;
mem[16'hCD27] = 8'h00;
mem[16'hCD28] = 8'h00;
mem[16'hCD29] = 8'h00;
mem[16'hCD2A] = 8'h00;
mem[16'hCD2B] = 8'h00;
mem[16'hCD2C] = 8'h00;
mem[16'hCD2D] = 8'h00;
mem[16'hCD2E] = 8'h00;
mem[16'hCD2F] = 8'h00;
mem[16'hCD30] = 8'h00;
mem[16'hCD31] = 8'h00;
mem[16'hCD32] = 8'h00;
mem[16'hCD33] = 8'h00;
mem[16'hCD34] = 8'h00;
mem[16'hCD35] = 8'h00;
mem[16'hCD36] = 8'h00;
mem[16'hCD37] = 8'h00;
mem[16'hCD38] = 8'h00;
mem[16'hCD39] = 8'h00;
mem[16'hCD3A] = 8'h00;
mem[16'hCD3B] = 8'h00;
mem[16'hCD3C] = 8'h00;
mem[16'hCD3D] = 8'h00;
mem[16'hCD3E] = 8'h00;
mem[16'hCD3F] = 8'h00;
mem[16'hCD40] = 8'h00;
mem[16'hCD41] = 8'h00;
mem[16'hCD42] = 8'h00;
mem[16'hCD43] = 8'h00;
mem[16'hCD44] = 8'h00;
mem[16'hCD45] = 8'h00;
mem[16'hCD46] = 8'h00;
mem[16'hCD47] = 8'h00;
mem[16'hCD48] = 8'h00;
mem[16'hCD49] = 8'h00;
mem[16'hCD4A] = 8'h00;
mem[16'hCD4B] = 8'h00;
mem[16'hCD4C] = 8'h00;
mem[16'hCD4D] = 8'h00;
mem[16'hCD4E] = 8'h00;
mem[16'hCD4F] = 8'h00;
mem[16'hCD50] = 8'h00;
mem[16'hCD51] = 8'h00;
mem[16'hCD52] = 8'h00;
mem[16'hCD53] = 8'h00;
mem[16'hCD54] = 8'h00;
mem[16'hCD55] = 8'h00;
mem[16'hCD56] = 8'h00;
mem[16'hCD57] = 8'h00;
mem[16'hCD58] = 8'h00;
mem[16'hCD59] = 8'h00;
mem[16'hCD5A] = 8'h00;
mem[16'hCD5B] = 8'h00;
mem[16'hCD5C] = 8'h00;
mem[16'hCD5D] = 8'h00;
mem[16'hCD5E] = 8'h00;
mem[16'hCD5F] = 8'h00;
mem[16'hCD60] = 8'h00;
mem[16'hCD61] = 8'h00;
mem[16'hCD62] = 8'h00;
mem[16'hCD63] = 8'h00;
mem[16'hCD64] = 8'h00;
mem[16'hCD65] = 8'h00;
mem[16'hCD66] = 8'h00;
mem[16'hCD67] = 8'h00;
mem[16'hCD68] = 8'h00;
mem[16'hCD69] = 8'h00;
mem[16'hCD6A] = 8'h00;
mem[16'hCD6B] = 8'h00;
mem[16'hCD6C] = 8'h00;
mem[16'hCD6D] = 8'h00;
mem[16'hCD6E] = 8'h00;
mem[16'hCD6F] = 8'h00;
mem[16'hCD70] = 8'h00;
mem[16'hCD71] = 8'h00;
mem[16'hCD72] = 8'h00;
mem[16'hCD73] = 8'h00;
mem[16'hCD74] = 8'h00;
mem[16'hCD75] = 8'h00;
mem[16'hCD76] = 8'h00;
mem[16'hCD77] = 8'h00;
mem[16'hCD78] = 8'h00;
mem[16'hCD79] = 8'h00;
mem[16'hCD7A] = 8'h00;
mem[16'hCD7B] = 8'h00;
mem[16'hCD7C] = 8'h00;
mem[16'hCD7D] = 8'h00;
mem[16'hCD7E] = 8'h00;
mem[16'hCD7F] = 8'h00;
mem[16'hCD80] = 8'h00;
mem[16'hCD81] = 8'h00;
mem[16'hCD82] = 8'h00;
mem[16'hCD83] = 8'h00;
mem[16'hCD84] = 8'h00;
mem[16'hCD85] = 8'h00;
mem[16'hCD86] = 8'h00;
mem[16'hCD87] = 8'h00;
mem[16'hCD88] = 8'h00;
mem[16'hCD89] = 8'h00;
mem[16'hCD8A] = 8'h00;
mem[16'hCD8B] = 8'h00;
mem[16'hCD8C] = 8'h00;
mem[16'hCD8D] = 8'h00;
mem[16'hCD8E] = 8'h00;
mem[16'hCD8F] = 8'h00;
mem[16'hCD90] = 8'h00;
mem[16'hCD91] = 8'h00;
mem[16'hCD92] = 8'h00;
mem[16'hCD93] = 8'h00;
mem[16'hCD94] = 8'h00;
mem[16'hCD95] = 8'h00;
mem[16'hCD96] = 8'h00;
mem[16'hCD97] = 8'h00;
mem[16'hCD98] = 8'h00;
mem[16'hCD99] = 8'h00;
mem[16'hCD9A] = 8'h00;
mem[16'hCD9B] = 8'h00;
mem[16'hCD9C] = 8'h00;
mem[16'hCD9D] = 8'h00;
mem[16'hCD9E] = 8'h00;
mem[16'hCD9F] = 8'h00;
mem[16'hCDA0] = 8'h00;
mem[16'hCDA1] = 8'h00;
mem[16'hCDA2] = 8'h00;
mem[16'hCDA3] = 8'h00;
mem[16'hCDA4] = 8'h00;
mem[16'hCDA5] = 8'h00;
mem[16'hCDA6] = 8'h00;
mem[16'hCDA7] = 8'h00;
mem[16'hCDA8] = 8'h00;
mem[16'hCDA9] = 8'h00;
mem[16'hCDAA] = 8'h00;
mem[16'hCDAB] = 8'h00;
mem[16'hCDAC] = 8'h00;
mem[16'hCDAD] = 8'h00;
mem[16'hCDAE] = 8'h00;
mem[16'hCDAF] = 8'h00;
mem[16'hCDB0] = 8'h00;
mem[16'hCDB1] = 8'h00;
mem[16'hCDB2] = 8'h00;
mem[16'hCDB3] = 8'h00;
mem[16'hCDB4] = 8'h00;
mem[16'hCDB5] = 8'h00;
mem[16'hCDB6] = 8'h00;
mem[16'hCDB7] = 8'h00;
mem[16'hCDB8] = 8'h00;
mem[16'hCDB9] = 8'h00;
mem[16'hCDBA] = 8'h00;
mem[16'hCDBB] = 8'h00;
mem[16'hCDBC] = 8'h00;
mem[16'hCDBD] = 8'h00;
mem[16'hCDBE] = 8'h00;
mem[16'hCDBF] = 8'h00;
mem[16'hCDC0] = 8'h00;
mem[16'hCDC1] = 8'h00;
mem[16'hCDC2] = 8'h00;
mem[16'hCDC3] = 8'h00;
mem[16'hCDC4] = 8'h00;
mem[16'hCDC5] = 8'h00;
mem[16'hCDC6] = 8'h00;
mem[16'hCDC7] = 8'h00;
mem[16'hCDC8] = 8'h00;
mem[16'hCDC9] = 8'h00;
mem[16'hCDCA] = 8'h00;
mem[16'hCDCB] = 8'h00;
mem[16'hCDCC] = 8'h00;
mem[16'hCDCD] = 8'h00;
mem[16'hCDCE] = 8'h00;
mem[16'hCDCF] = 8'h00;
mem[16'hCDD0] = 8'h00;
mem[16'hCDD1] = 8'h00;
mem[16'hCDD2] = 8'h00;
mem[16'hCDD3] = 8'h00;
mem[16'hCDD4] = 8'h00;
mem[16'hCDD5] = 8'h00;
mem[16'hCDD6] = 8'h00;
mem[16'hCDD7] = 8'h00;
mem[16'hCDD8] = 8'h00;
mem[16'hCDD9] = 8'h00;
mem[16'hCDDA] = 8'h00;
mem[16'hCDDB] = 8'h00;
mem[16'hCDDC] = 8'h00;
mem[16'hCDDD] = 8'h00;
mem[16'hCDDE] = 8'h00;
mem[16'hCDDF] = 8'h00;
mem[16'hCDE0] = 8'h00;
mem[16'hCDE1] = 8'h00;
mem[16'hCDE2] = 8'h00;
mem[16'hCDE3] = 8'h00;
mem[16'hCDE4] = 8'h00;
mem[16'hCDE5] = 8'h00;
mem[16'hCDE6] = 8'h00;
mem[16'hCDE7] = 8'h00;
mem[16'hCDE8] = 8'h00;
mem[16'hCDE9] = 8'h00;
mem[16'hCDEA] = 8'h00;
mem[16'hCDEB] = 8'h00;
mem[16'hCDEC] = 8'h00;
mem[16'hCDED] = 8'h00;
mem[16'hCDEE] = 8'h00;
mem[16'hCDEF] = 8'h00;
mem[16'hCDF0] = 8'h00;
mem[16'hCDF1] = 8'h00;
mem[16'hCDF2] = 8'h00;
mem[16'hCDF3] = 8'h00;
mem[16'hCDF4] = 8'h00;
mem[16'hCDF5] = 8'h00;
mem[16'hCDF6] = 8'h00;
mem[16'hCDF7] = 8'h00;
mem[16'hCDF8] = 8'h00;
mem[16'hCDF9] = 8'h00;
mem[16'hCDFA] = 8'h00;
mem[16'hCDFB] = 8'h00;
mem[16'hCDFC] = 8'h00;
mem[16'hCDFD] = 8'h00;
mem[16'hCDFE] = 8'h00;
mem[16'hCDFF] = 8'h00;
mem[16'hCE00] = 8'h00;
mem[16'hCE01] = 8'h00;
mem[16'hCE02] = 8'h00;
mem[16'hCE03] = 8'h00;
mem[16'hCE04] = 8'h00;
mem[16'hCE05] = 8'h00;
mem[16'hCE06] = 8'h00;
mem[16'hCE07] = 8'h00;
mem[16'hCE08] = 8'h00;
mem[16'hCE09] = 8'h00;
mem[16'hCE0A] = 8'h00;
mem[16'hCE0B] = 8'h00;
mem[16'hCE0C] = 8'h00;
mem[16'hCE0D] = 8'h00;
mem[16'hCE0E] = 8'h00;
mem[16'hCE0F] = 8'h00;
mem[16'hCE10] = 8'h00;
mem[16'hCE11] = 8'h00;
mem[16'hCE12] = 8'h00;
mem[16'hCE13] = 8'h00;
mem[16'hCE14] = 8'h00;
mem[16'hCE15] = 8'h00;
mem[16'hCE16] = 8'h00;
mem[16'hCE17] = 8'h00;
mem[16'hCE18] = 8'h00;
mem[16'hCE19] = 8'h00;
mem[16'hCE1A] = 8'h00;
mem[16'hCE1B] = 8'h00;
mem[16'hCE1C] = 8'h00;
mem[16'hCE1D] = 8'h00;
mem[16'hCE1E] = 8'h00;
mem[16'hCE1F] = 8'h00;
mem[16'hCE20] = 8'h00;
mem[16'hCE21] = 8'h00;
mem[16'hCE22] = 8'h00;
mem[16'hCE23] = 8'h00;
mem[16'hCE24] = 8'h00;
mem[16'hCE25] = 8'h00;
mem[16'hCE26] = 8'h00;
mem[16'hCE27] = 8'h00;
mem[16'hCE28] = 8'h00;
mem[16'hCE29] = 8'h00;
mem[16'hCE2A] = 8'h00;
mem[16'hCE2B] = 8'h00;
mem[16'hCE2C] = 8'h00;
mem[16'hCE2D] = 8'h00;
mem[16'hCE2E] = 8'h00;
mem[16'hCE2F] = 8'h00;
mem[16'hCE30] = 8'h00;
mem[16'hCE31] = 8'h00;
mem[16'hCE32] = 8'h00;
mem[16'hCE33] = 8'h00;
mem[16'hCE34] = 8'h00;
mem[16'hCE35] = 8'h00;
mem[16'hCE36] = 8'h00;
mem[16'hCE37] = 8'h00;
mem[16'hCE38] = 8'h00;
mem[16'hCE39] = 8'h00;
mem[16'hCE3A] = 8'h00;
mem[16'hCE3B] = 8'h00;
mem[16'hCE3C] = 8'h00;
mem[16'hCE3D] = 8'h00;
mem[16'hCE3E] = 8'h00;
mem[16'hCE3F] = 8'h00;
mem[16'hCE40] = 8'h00;
mem[16'hCE41] = 8'h00;
mem[16'hCE42] = 8'h00;
mem[16'hCE43] = 8'h00;
mem[16'hCE44] = 8'h00;
mem[16'hCE45] = 8'h00;
mem[16'hCE46] = 8'h00;
mem[16'hCE47] = 8'h00;
mem[16'hCE48] = 8'h00;
mem[16'hCE49] = 8'h00;
mem[16'hCE4A] = 8'h00;
mem[16'hCE4B] = 8'h00;
mem[16'hCE4C] = 8'h00;
mem[16'hCE4D] = 8'h00;
mem[16'hCE4E] = 8'h00;
mem[16'hCE4F] = 8'h00;
mem[16'hCE50] = 8'h00;
mem[16'hCE51] = 8'h00;
mem[16'hCE52] = 8'h00;
mem[16'hCE53] = 8'h00;
mem[16'hCE54] = 8'h00;
mem[16'hCE55] = 8'h00;
mem[16'hCE56] = 8'h00;
mem[16'hCE57] = 8'h00;
mem[16'hCE58] = 8'h00;
mem[16'hCE59] = 8'h00;
mem[16'hCE5A] = 8'h00;
mem[16'hCE5B] = 8'h00;
mem[16'hCE5C] = 8'h00;
mem[16'hCE5D] = 8'h00;
mem[16'hCE5E] = 8'h00;
mem[16'hCE5F] = 8'h00;
mem[16'hCE60] = 8'h00;
mem[16'hCE61] = 8'h00;
mem[16'hCE62] = 8'h00;
mem[16'hCE63] = 8'h00;
mem[16'hCE64] = 8'h00;
mem[16'hCE65] = 8'h00;
mem[16'hCE66] = 8'h00;
mem[16'hCE67] = 8'h00;
mem[16'hCE68] = 8'h00;
mem[16'hCE69] = 8'h00;
mem[16'hCE6A] = 8'h00;
mem[16'hCE6B] = 8'h00;
mem[16'hCE6C] = 8'h00;
mem[16'hCE6D] = 8'h00;
mem[16'hCE6E] = 8'h00;
mem[16'hCE6F] = 8'h00;
mem[16'hCE70] = 8'h00;
mem[16'hCE71] = 8'h00;
mem[16'hCE72] = 8'h00;
mem[16'hCE73] = 8'h00;
mem[16'hCE74] = 8'h00;
mem[16'hCE75] = 8'h00;
mem[16'hCE76] = 8'h00;
mem[16'hCE77] = 8'h00;
mem[16'hCE78] = 8'h00;
mem[16'hCE79] = 8'h00;
mem[16'hCE7A] = 8'h00;
mem[16'hCE7B] = 8'h00;
mem[16'hCE7C] = 8'h00;
mem[16'hCE7D] = 8'h00;
mem[16'hCE7E] = 8'h00;
mem[16'hCE7F] = 8'h00;
mem[16'hCE80] = 8'h00;
mem[16'hCE81] = 8'h00;
mem[16'hCE82] = 8'h00;
mem[16'hCE83] = 8'h00;
mem[16'hCE84] = 8'h00;
mem[16'hCE85] = 8'h00;
mem[16'hCE86] = 8'h00;
mem[16'hCE87] = 8'h00;
mem[16'hCE88] = 8'h00;
mem[16'hCE89] = 8'h00;
mem[16'hCE8A] = 8'h00;
mem[16'hCE8B] = 8'h00;
mem[16'hCE8C] = 8'h00;
mem[16'hCE8D] = 8'h00;
mem[16'hCE8E] = 8'h00;
mem[16'hCE8F] = 8'h00;
mem[16'hCE90] = 8'h00;
mem[16'hCE91] = 8'h00;
mem[16'hCE92] = 8'h00;
mem[16'hCE93] = 8'h00;
mem[16'hCE94] = 8'h00;
mem[16'hCE95] = 8'h00;
mem[16'hCE96] = 8'h00;
mem[16'hCE97] = 8'h00;
mem[16'hCE98] = 8'h00;
mem[16'hCE99] = 8'h00;
mem[16'hCE9A] = 8'h00;
mem[16'hCE9B] = 8'h00;
mem[16'hCE9C] = 8'h00;
mem[16'hCE9D] = 8'h00;
mem[16'hCE9E] = 8'h00;
mem[16'hCE9F] = 8'h00;
mem[16'hCEA0] = 8'h00;
mem[16'hCEA1] = 8'h00;
mem[16'hCEA2] = 8'h00;
mem[16'hCEA3] = 8'h00;
mem[16'hCEA4] = 8'h00;
mem[16'hCEA5] = 8'h00;
mem[16'hCEA6] = 8'h00;
mem[16'hCEA7] = 8'h00;
mem[16'hCEA8] = 8'h00;
mem[16'hCEA9] = 8'h00;
mem[16'hCEAA] = 8'h00;
mem[16'hCEAB] = 8'h00;
mem[16'hCEAC] = 8'h00;
mem[16'hCEAD] = 8'h00;
mem[16'hCEAE] = 8'h00;
mem[16'hCEAF] = 8'h00;
mem[16'hCEB0] = 8'h00;
mem[16'hCEB1] = 8'h00;
mem[16'hCEB2] = 8'h00;
mem[16'hCEB3] = 8'h00;
mem[16'hCEB4] = 8'h00;
mem[16'hCEB5] = 8'h00;
mem[16'hCEB6] = 8'h00;
mem[16'hCEB7] = 8'h00;
mem[16'hCEB8] = 8'h00;
mem[16'hCEB9] = 8'h00;
mem[16'hCEBA] = 8'h00;
mem[16'hCEBB] = 8'h00;
mem[16'hCEBC] = 8'h00;
mem[16'hCEBD] = 8'h00;
mem[16'hCEBE] = 8'h00;
mem[16'hCEBF] = 8'h00;
mem[16'hCEC0] = 8'h00;
mem[16'hCEC1] = 8'h00;
mem[16'hCEC2] = 8'h00;
mem[16'hCEC3] = 8'h00;
mem[16'hCEC4] = 8'h00;
mem[16'hCEC5] = 8'h00;
mem[16'hCEC6] = 8'h00;
mem[16'hCEC7] = 8'h00;
mem[16'hCEC8] = 8'h00;
mem[16'hCEC9] = 8'h00;
mem[16'hCECA] = 8'h00;
mem[16'hCECB] = 8'h00;
mem[16'hCECC] = 8'h00;
mem[16'hCECD] = 8'h00;
mem[16'hCECE] = 8'h00;
mem[16'hCECF] = 8'h00;
mem[16'hCED0] = 8'h00;
mem[16'hCED1] = 8'h00;
mem[16'hCED2] = 8'h00;
mem[16'hCED3] = 8'h00;
mem[16'hCED4] = 8'h00;
mem[16'hCED5] = 8'h00;
mem[16'hCED6] = 8'h00;
mem[16'hCED7] = 8'h00;
mem[16'hCED8] = 8'h00;
mem[16'hCED9] = 8'h00;
mem[16'hCEDA] = 8'h00;
mem[16'hCEDB] = 8'h00;
mem[16'hCEDC] = 8'h00;
mem[16'hCEDD] = 8'h00;
mem[16'hCEDE] = 8'h00;
mem[16'hCEDF] = 8'h00;
mem[16'hCEE0] = 8'h00;
mem[16'hCEE1] = 8'h00;
mem[16'hCEE2] = 8'h00;
mem[16'hCEE3] = 8'h00;
mem[16'hCEE4] = 8'h00;
mem[16'hCEE5] = 8'h00;
mem[16'hCEE6] = 8'h00;
mem[16'hCEE7] = 8'h00;
mem[16'hCEE8] = 8'h00;
mem[16'hCEE9] = 8'h00;
mem[16'hCEEA] = 8'h00;
mem[16'hCEEB] = 8'h00;
mem[16'hCEEC] = 8'h00;
mem[16'hCEED] = 8'h00;
mem[16'hCEEE] = 8'h00;
mem[16'hCEEF] = 8'h00;
mem[16'hCEF0] = 8'h00;
mem[16'hCEF1] = 8'h00;
mem[16'hCEF2] = 8'h00;
mem[16'hCEF3] = 8'h00;
mem[16'hCEF4] = 8'h00;
mem[16'hCEF5] = 8'h00;
mem[16'hCEF6] = 8'h00;
mem[16'hCEF7] = 8'h00;
mem[16'hCEF8] = 8'h00;
mem[16'hCEF9] = 8'h00;
mem[16'hCEFA] = 8'h00;
mem[16'hCEFB] = 8'h00;
mem[16'hCEFC] = 8'h00;
mem[16'hCEFD] = 8'h00;
mem[16'hCEFE] = 8'h00;
mem[16'hCEFF] = 8'h00;
mem[16'hCF00] = 8'h00;
mem[16'hCF01] = 8'h00;
mem[16'hCF02] = 8'h00;
mem[16'hCF03] = 8'h00;
mem[16'hCF04] = 8'h00;
mem[16'hCF05] = 8'h00;
mem[16'hCF06] = 8'h00;
mem[16'hCF07] = 8'h00;
mem[16'hCF08] = 8'h00;
mem[16'hCF09] = 8'h00;
mem[16'hCF0A] = 8'h00;
mem[16'hCF0B] = 8'h00;
mem[16'hCF0C] = 8'h00;
mem[16'hCF0D] = 8'h00;
mem[16'hCF0E] = 8'h00;
mem[16'hCF0F] = 8'h00;
mem[16'hCF10] = 8'h00;
mem[16'hCF11] = 8'h00;
mem[16'hCF12] = 8'h00;
mem[16'hCF13] = 8'h00;
mem[16'hCF14] = 8'h00;
mem[16'hCF15] = 8'h00;
mem[16'hCF16] = 8'h00;
mem[16'hCF17] = 8'h00;
mem[16'hCF18] = 8'h00;
mem[16'hCF19] = 8'h00;
mem[16'hCF1A] = 8'h00;
mem[16'hCF1B] = 8'h00;
mem[16'hCF1C] = 8'h00;
mem[16'hCF1D] = 8'h00;
mem[16'hCF1E] = 8'h00;
mem[16'hCF1F] = 8'h00;
mem[16'hCF20] = 8'h00;
mem[16'hCF21] = 8'h00;
mem[16'hCF22] = 8'h00;
mem[16'hCF23] = 8'h00;
mem[16'hCF24] = 8'h00;
mem[16'hCF25] = 8'h00;
mem[16'hCF26] = 8'h00;
mem[16'hCF27] = 8'h00;
mem[16'hCF28] = 8'h00;
mem[16'hCF29] = 8'h00;
mem[16'hCF2A] = 8'h00;
mem[16'hCF2B] = 8'h00;
mem[16'hCF2C] = 8'h00;
mem[16'hCF2D] = 8'h00;
mem[16'hCF2E] = 8'h00;
mem[16'hCF2F] = 8'h00;
mem[16'hCF30] = 8'h00;
mem[16'hCF31] = 8'h00;
mem[16'hCF32] = 8'h00;
mem[16'hCF33] = 8'h00;
mem[16'hCF34] = 8'h00;
mem[16'hCF35] = 8'h00;
mem[16'hCF36] = 8'h00;
mem[16'hCF37] = 8'h00;
mem[16'hCF38] = 8'h00;
mem[16'hCF39] = 8'h00;
mem[16'hCF3A] = 8'h00;
mem[16'hCF3B] = 8'h00;
mem[16'hCF3C] = 8'h00;
mem[16'hCF3D] = 8'h00;
mem[16'hCF3E] = 8'h00;
mem[16'hCF3F] = 8'h00;
mem[16'hCF40] = 8'h00;
mem[16'hCF41] = 8'h00;
mem[16'hCF42] = 8'h00;
mem[16'hCF43] = 8'h00;
mem[16'hCF44] = 8'h00;
mem[16'hCF45] = 8'h00;
mem[16'hCF46] = 8'h00;
mem[16'hCF47] = 8'h00;
mem[16'hCF48] = 8'h00;
mem[16'hCF49] = 8'h00;
mem[16'hCF4A] = 8'h00;
mem[16'hCF4B] = 8'h00;
mem[16'hCF4C] = 8'h00;
mem[16'hCF4D] = 8'h00;
mem[16'hCF4E] = 8'h00;
mem[16'hCF4F] = 8'h00;
mem[16'hCF50] = 8'h00;
mem[16'hCF51] = 8'h00;
mem[16'hCF52] = 8'h00;
mem[16'hCF53] = 8'h00;
mem[16'hCF54] = 8'h00;
mem[16'hCF55] = 8'h00;
mem[16'hCF56] = 8'h00;
mem[16'hCF57] = 8'h00;
mem[16'hCF58] = 8'h00;
mem[16'hCF59] = 8'h00;
mem[16'hCF5A] = 8'h00;
mem[16'hCF5B] = 8'h00;
mem[16'hCF5C] = 8'h00;
mem[16'hCF5D] = 8'h00;
mem[16'hCF5E] = 8'h00;
mem[16'hCF5F] = 8'h00;
mem[16'hCF60] = 8'h00;
mem[16'hCF61] = 8'h00;
mem[16'hCF62] = 8'h00;
mem[16'hCF63] = 8'h00;
mem[16'hCF64] = 8'h00;
mem[16'hCF65] = 8'h00;
mem[16'hCF66] = 8'h00;
mem[16'hCF67] = 8'h00;
mem[16'hCF68] = 8'h00;
mem[16'hCF69] = 8'h00;
mem[16'hCF6A] = 8'h00;
mem[16'hCF6B] = 8'h00;
mem[16'hCF6C] = 8'h00;
mem[16'hCF6D] = 8'h00;
mem[16'hCF6E] = 8'h00;
mem[16'hCF6F] = 8'h00;
mem[16'hCF70] = 8'h00;
mem[16'hCF71] = 8'h00;
mem[16'hCF72] = 8'h00;
mem[16'hCF73] = 8'h00;
mem[16'hCF74] = 8'h00;
mem[16'hCF75] = 8'h00;
mem[16'hCF76] = 8'h00;
mem[16'hCF77] = 8'h00;
mem[16'hCF78] = 8'h00;
mem[16'hCF79] = 8'h00;
mem[16'hCF7A] = 8'h00;
mem[16'hCF7B] = 8'h00;
mem[16'hCF7C] = 8'h00;
mem[16'hCF7D] = 8'h00;
mem[16'hCF7E] = 8'h00;
mem[16'hCF7F] = 8'h00;
mem[16'hCF80] = 8'h00;
mem[16'hCF81] = 8'h00;
mem[16'hCF82] = 8'h00;
mem[16'hCF83] = 8'h00;
mem[16'hCF84] = 8'h00;
mem[16'hCF85] = 8'h00;
mem[16'hCF86] = 8'h00;
mem[16'hCF87] = 8'h00;
mem[16'hCF88] = 8'h00;
mem[16'hCF89] = 8'h00;
mem[16'hCF8A] = 8'h00;
mem[16'hCF8B] = 8'h00;
mem[16'hCF8C] = 8'h00;
mem[16'hCF8D] = 8'h00;
mem[16'hCF8E] = 8'h00;
mem[16'hCF8F] = 8'h00;
mem[16'hCF90] = 8'h00;
mem[16'hCF91] = 8'h00;
mem[16'hCF92] = 8'h00;
mem[16'hCF93] = 8'h00;
mem[16'hCF94] = 8'h00;
mem[16'hCF95] = 8'h00;
mem[16'hCF96] = 8'h00;
mem[16'hCF97] = 8'h00;
mem[16'hCF98] = 8'h00;
mem[16'hCF99] = 8'h00;
mem[16'hCF9A] = 8'h00;
mem[16'hCF9B] = 8'h00;
mem[16'hCF9C] = 8'h00;
mem[16'hCF9D] = 8'h00;
mem[16'hCF9E] = 8'h00;
mem[16'hCF9F] = 8'h00;
mem[16'hCFA0] = 8'h00;
mem[16'hCFA1] = 8'h00;
mem[16'hCFA2] = 8'h00;
mem[16'hCFA3] = 8'h00;
mem[16'hCFA4] = 8'h00;
mem[16'hCFA5] = 8'h00;
mem[16'hCFA6] = 8'h00;
mem[16'hCFA7] = 8'h00;
mem[16'hCFA8] = 8'h00;
mem[16'hCFA9] = 8'h00;
mem[16'hCFAA] = 8'h00;
mem[16'hCFAB] = 8'h00;
mem[16'hCFAC] = 8'h00;
mem[16'hCFAD] = 8'h00;
mem[16'hCFAE] = 8'h00;
mem[16'hCFAF] = 8'h00;
mem[16'hCFB0] = 8'h00;
mem[16'hCFB1] = 8'h00;
mem[16'hCFB2] = 8'h00;
mem[16'hCFB3] = 8'h00;
mem[16'hCFB4] = 8'h00;
mem[16'hCFB5] = 8'h00;
mem[16'hCFB6] = 8'h00;
mem[16'hCFB7] = 8'h00;
mem[16'hCFB8] = 8'h00;
mem[16'hCFB9] = 8'h00;
mem[16'hCFBA] = 8'h00;
mem[16'hCFBB] = 8'h00;
mem[16'hCFBC] = 8'h00;
mem[16'hCFBD] = 8'h00;
mem[16'hCFBE] = 8'h00;
mem[16'hCFBF] = 8'h00;
mem[16'hCFC0] = 8'h00;
mem[16'hCFC1] = 8'h00;
mem[16'hCFC2] = 8'h00;
mem[16'hCFC3] = 8'h00;
mem[16'hCFC4] = 8'h00;
mem[16'hCFC5] = 8'h00;
mem[16'hCFC6] = 8'h00;
mem[16'hCFC7] = 8'h00;
mem[16'hCFC8] = 8'h00;
mem[16'hCFC9] = 8'h00;
mem[16'hCFCA] = 8'h00;
mem[16'hCFCB] = 8'h00;
mem[16'hCFCC] = 8'h00;
mem[16'hCFCD] = 8'h00;
mem[16'hCFCE] = 8'h00;
mem[16'hCFCF] = 8'h00;
mem[16'hCFD0] = 8'h00;
mem[16'hCFD1] = 8'h00;
mem[16'hCFD2] = 8'h00;
mem[16'hCFD3] = 8'h00;
mem[16'hCFD4] = 8'h00;
mem[16'hCFD5] = 8'h00;
mem[16'hCFD6] = 8'h00;
mem[16'hCFD7] = 8'h00;
mem[16'hCFD8] = 8'h00;
mem[16'hCFD9] = 8'h00;
mem[16'hCFDA] = 8'h00;
mem[16'hCFDB] = 8'h00;
mem[16'hCFDC] = 8'h00;
mem[16'hCFDD] = 8'h00;
mem[16'hCFDE] = 8'h00;
mem[16'hCFDF] = 8'h00;
mem[16'hCFE0] = 8'h00;
mem[16'hCFE1] = 8'h00;
mem[16'hCFE2] = 8'h00;
mem[16'hCFE3] = 8'h00;
mem[16'hCFE4] = 8'h00;
mem[16'hCFE5] = 8'h00;
mem[16'hCFE6] = 8'h00;
mem[16'hCFE7] = 8'h00;
mem[16'hCFE8] = 8'h00;
mem[16'hCFE9] = 8'h00;
mem[16'hCFEA] = 8'h00;
mem[16'hCFEB] = 8'h00;
mem[16'hCFEC] = 8'h00;
mem[16'hCFED] = 8'h00;
mem[16'hCFEE] = 8'h00;
mem[16'hCFEF] = 8'h00;
mem[16'hCFF0] = 8'h00;
mem[16'hCFF1] = 8'h00;
mem[16'hCFF2] = 8'h00;
mem[16'hCFF3] = 8'h00;
mem[16'hCFF4] = 8'h00;
mem[16'hCFF5] = 8'h00;
mem[16'hCFF6] = 8'h00;
mem[16'hCFF7] = 8'h00;
mem[16'hCFF8] = 8'h00;
mem[16'hCFF9] = 8'h00;
mem[16'hCFFA] = 8'h00;
mem[16'hCFFB] = 8'h00;
mem[16'hCFFC] = 8'h00;
mem[16'hCFFD] = 8'h00;
mem[16'hCFFE] = 8'h00;
mem[16'hCFFF] = 8'h00;
mem[16'hD000] = 8'h6F;
mem[16'hD001] = 8'hD8;
mem[16'hD002] = 8'h65;
mem[16'hD003] = 8'hD7;
mem[16'hD004] = 8'hF8;
mem[16'hD005] = 8'hDC;
mem[16'hD006] = 8'h94;
mem[16'hD007] = 8'hD9;
mem[16'hD008] = 8'hB1;
mem[16'hD009] = 8'hDB;
mem[16'hD00A] = 8'h30;
mem[16'hD00B] = 8'hF3;
mem[16'hD00C] = 8'hD8;
mem[16'hD00D] = 8'hDF;
mem[16'hD00E] = 8'hE1;
mem[16'hD00F] = 8'hDB;
mem[16'hD010] = 8'h8F;
mem[16'hD011] = 8'hF3;
mem[16'hD012] = 8'h98;
mem[16'hD013] = 8'hF3;
mem[16'hD014] = 8'hE4;
mem[16'hD015] = 8'hF1;
mem[16'hD016] = 8'hDD;
mem[16'hD017] = 8'hF1;
mem[16'hD018] = 8'hD4;
mem[16'hD019] = 8'hF1;
mem[16'hD01A] = 8'h24;
mem[16'hD01B] = 8'hF2;
mem[16'hD01C] = 8'h31;
mem[16'hD01D] = 8'hF2;
mem[16'hD01E] = 8'h40;
mem[16'hD01F] = 8'hF2;
mem[16'hD020] = 8'hD7;
mem[16'hD021] = 8'hF3;
mem[16'hD022] = 8'hE1;
mem[16'hD023] = 8'hF3;
mem[16'hD024] = 8'hE8;
mem[16'hD025] = 8'hF6;
mem[16'hD026] = 8'hFD;
mem[16'hD027] = 8'hF6;
mem[16'hD028] = 8'h68;
mem[16'hD029] = 8'hF7;
mem[16'hD02A] = 8'h6E;
mem[16'hD02B] = 8'hF7;
mem[16'hD02C] = 8'hE6;
mem[16'hD02D] = 8'hF7;
mem[16'hD02E] = 8'h57;
mem[16'hD02F] = 8'hFC;
mem[16'hD030] = 8'h20;
mem[16'hD031] = 8'hF7;
mem[16'hD032] = 8'h26;
mem[16'hD033] = 8'hF7;
mem[16'hD034] = 8'h74;
mem[16'hD035] = 8'hF7;
mem[16'hD036] = 8'h6C;
mem[16'hD037] = 8'hF2;
mem[16'hD038] = 8'h6E;
mem[16'hD039] = 8'hF2;
mem[16'hD03A] = 8'h72;
mem[16'hD03B] = 8'hF2;
mem[16'hD03C] = 8'h76;
mem[16'hD03D] = 8'hF2;
mem[16'hD03E] = 8'h7F;
mem[16'hD03F] = 8'hF2;
mem[16'hD040] = 8'h4E;
mem[16'hD041] = 8'hF2;
mem[16'hD042] = 8'h6A;
mem[16'hD043] = 8'hD9;
mem[16'hD044] = 8'h55;
mem[16'hD045] = 8'hF2;
mem[16'hD046] = 8'h85;
mem[16'hD047] = 8'hF2;
mem[16'hD048] = 8'hA5;
mem[16'hD049] = 8'hF2;
mem[16'hD04A] = 8'hCA;
mem[16'hD04B] = 8'hF2;
mem[16'hD04C] = 8'h17;
mem[16'hD04D] = 8'hF3;
mem[16'hD04E] = 8'hBB;
mem[16'hD04F] = 8'hF3;
mem[16'hD050] = 8'h9E;
mem[16'hD051] = 8'hF3;
mem[16'hD052] = 8'h61;
mem[16'hD053] = 8'hF2;
mem[16'hD054] = 8'h45;
mem[16'hD055] = 8'hDA;
mem[16'hD056] = 8'h3D;
mem[16'hD057] = 8'hD9;
mem[16'hD058] = 8'h11;
mem[16'hD059] = 8'hD9;
mem[16'hD05A] = 8'hC8;
mem[16'hD05B] = 8'hD9;
mem[16'hD05C] = 8'h48;
mem[16'hD05D] = 8'hD8;
mem[16'hD05E] = 8'hF4;
mem[16'hD05F] = 8'h03;
mem[16'hD060] = 8'h20;
mem[16'hD061] = 8'hD9;
mem[16'hD062] = 8'h6A;
mem[16'hD063] = 8'hD9;
mem[16'hD064] = 8'hDB;
mem[16'hD065] = 8'hD9;
mem[16'hD066] = 8'h6D;
mem[16'hD067] = 8'hD8;
mem[16'hD068] = 8'hEB;
mem[16'hD069] = 8'hD9;
mem[16'hD06A] = 8'h83;
mem[16'hD06B] = 8'hE7;
mem[16'hD06C] = 8'hC8;
mem[16'hD06D] = 8'hD8;
mem[16'hD06E] = 8'hAF;
mem[16'hD06F] = 8'hD8;
mem[16'hD070] = 8'h12;
mem[16'hD071] = 8'hE3;
mem[16'hD072] = 8'h7A;
mem[16'hD073] = 8'hE7;
mem[16'hD074] = 8'hD4;
mem[16'hD075] = 8'hDA;
mem[16'hD076] = 8'h95;
mem[16'hD077] = 8'hD8;
mem[16'hD078] = 8'hA4;
mem[16'hD079] = 8'hD6;
mem[16'hD07A] = 8'h69;
mem[16'hD07B] = 8'hD6;
mem[16'hD07C] = 8'h9F;
mem[16'hD07D] = 8'hDB;
mem[16'hD07E] = 8'h48;
mem[16'hD07F] = 8'hD6;
mem[16'hD080] = 8'h90;
mem[16'hD081] = 8'hEB;
mem[16'hD082] = 8'h23;
mem[16'hD083] = 8'hEC;
mem[16'hD084] = 8'hAF;
mem[16'hD085] = 8'hEB;
mem[16'hD086] = 8'h0A;
mem[16'hD087] = 8'h00;
mem[16'hD088] = 8'hDE;
mem[16'hD089] = 8'hE2;
mem[16'hD08A] = 8'h12;
mem[16'hD08B] = 8'hD4;
mem[16'hD08C] = 8'hCD;
mem[16'hD08D] = 8'hDF;
mem[16'hD08E] = 8'hFF;
mem[16'hD08F] = 8'hE2;
mem[16'hD090] = 8'h8D;
mem[16'hD091] = 8'hEE;
mem[16'hD092] = 8'hAE;
mem[16'hD093] = 8'hEF;
mem[16'hD094] = 8'h41;
mem[16'hD095] = 8'hE9;
mem[16'hD096] = 8'h09;
mem[16'hD097] = 8'hEF;
mem[16'hD098] = 8'hEA;
mem[16'hD099] = 8'hEF;
mem[16'hD09A] = 8'hF1;
mem[16'hD09B] = 8'hEF;
mem[16'hD09C] = 8'h3A;
mem[16'hD09D] = 8'hF0;
mem[16'hD09E] = 8'h9E;
mem[16'hD09F] = 8'hF0;
mem[16'hD0A0] = 8'h64;
mem[16'hD0A1] = 8'hE7;
mem[16'hD0A2] = 8'hD6;
mem[16'hD0A3] = 8'hE6;
mem[16'hD0A4] = 8'hC5;
mem[16'hD0A5] = 8'hE3;
mem[16'hD0A6] = 8'h07;
mem[16'hD0A7] = 8'hE7;
mem[16'hD0A8] = 8'hE5;
mem[16'hD0A9] = 8'hE6;
mem[16'hD0AA] = 8'h46;
mem[16'hD0AB] = 8'hE6;
mem[16'hD0AC] = 8'h5A;
mem[16'hD0AD] = 8'hE6;
mem[16'hD0AE] = 8'h86;
mem[16'hD0AF] = 8'hE6;
mem[16'hD0B0] = 8'h91;
mem[16'hD0B1] = 8'hE6;
mem[16'hD0B2] = 8'h79;
mem[16'hD0B3] = 8'hC0;
mem[16'hD0B4] = 8'hE7;
mem[16'hD0B5] = 8'h79;
mem[16'hD0B6] = 8'hA9;
mem[16'hD0B7] = 8'hE7;
mem[16'hD0B8] = 8'h7B;
mem[16'hD0B9] = 8'h81;
mem[16'hD0BA] = 8'hE9;
mem[16'hD0BB] = 8'h7B;
mem[16'hD0BC] = 8'h68;
mem[16'hD0BD] = 8'hEA;
mem[16'hD0BE] = 8'h7D;
mem[16'hD0BF] = 8'h96;
mem[16'hD0C0] = 8'hEE;
mem[16'hD0C1] = 8'h50;
mem[16'hD0C2] = 8'h54;
mem[16'hD0C3] = 8'hDF;
mem[16'hD0C4] = 8'h46;
mem[16'hD0C5] = 8'h4E;
mem[16'hD0C6] = 8'hDF;
mem[16'hD0C7] = 8'h7F;
mem[16'hD0C8] = 8'hCF;
mem[16'hD0C9] = 8'hEE;
mem[16'hD0CA] = 8'h7F;
mem[16'hD0CB] = 8'h97;
mem[16'hD0CC] = 8'hDE;
mem[16'hD0CD] = 8'h64;
mem[16'hD0CE] = 8'h64;
mem[16'hD0CF] = 8'hDF;
mem[16'hD0D0] = 8'h45;
mem[16'hD0D1] = 8'h4E;
mem[16'hD0D2] = 8'hC4;
mem[16'hD0D3] = 8'h46;
mem[16'hD0D4] = 8'h4F;
mem[16'hD0D5] = 8'hD2;
mem[16'hD0D6] = 8'h4E;
mem[16'hD0D7] = 8'h45;
mem[16'hD0D8] = 8'h58;
mem[16'hD0D9] = 8'hD4;
mem[16'hD0DA] = 8'h44;
mem[16'hD0DB] = 8'h41;
mem[16'hD0DC] = 8'h54;
mem[16'hD0DD] = 8'hC1;
mem[16'hD0DE] = 8'h49;
mem[16'hD0DF] = 8'h4E;
mem[16'hD0E0] = 8'h50;
mem[16'hD0E1] = 8'h55;
mem[16'hD0E2] = 8'hD4;
mem[16'hD0E3] = 8'h44;
mem[16'hD0E4] = 8'h45;
mem[16'hD0E5] = 8'hCC;
mem[16'hD0E6] = 8'h44;
mem[16'hD0E7] = 8'h49;
mem[16'hD0E8] = 8'hCD;
mem[16'hD0E9] = 8'h52;
mem[16'hD0EA] = 8'h45;
mem[16'hD0EB] = 8'h41;
mem[16'hD0EC] = 8'hC4;
mem[16'hD0ED] = 8'h47;
mem[16'hD0EE] = 8'hD2;
mem[16'hD0EF] = 8'h54;
mem[16'hD0F0] = 8'h45;
mem[16'hD0F1] = 8'h58;
mem[16'hD0F2] = 8'hD4;
mem[16'hD0F3] = 8'h50;
mem[16'hD0F4] = 8'h52;
mem[16'hD0F5] = 8'hA3;
mem[16'hD0F6] = 8'h49;
mem[16'hD0F7] = 8'h4E;
mem[16'hD0F8] = 8'hA3;
mem[16'hD0F9] = 8'h43;
mem[16'hD0FA] = 8'h41;
mem[16'hD0FB] = 8'h4C;
mem[16'hD0FC] = 8'hCC;
mem[16'hD0FD] = 8'h50;
mem[16'hD0FE] = 8'h4C;
mem[16'hD0FF] = 8'h4F;
mem[16'hD100] = 8'hD4;
mem[16'hD101] = 8'h48;
mem[16'hD102] = 8'h4C;
mem[16'hD103] = 8'h49;
mem[16'hD104] = 8'hCE;
mem[16'hD105] = 8'h56;
mem[16'hD106] = 8'h4C;
mem[16'hD107] = 8'h49;
mem[16'hD108] = 8'hCE;
mem[16'hD109] = 8'h48;
mem[16'hD10A] = 8'h47;
mem[16'hD10B] = 8'h52;
mem[16'hD10C] = 8'hB2;
mem[16'hD10D] = 8'h48;
mem[16'hD10E] = 8'h47;
mem[16'hD10F] = 8'hD2;
mem[16'hD110] = 8'h48;
mem[16'hD111] = 8'h43;
mem[16'hD112] = 8'h4F;
mem[16'hD113] = 8'h4C;
mem[16'hD114] = 8'h4F;
mem[16'hD115] = 8'h52;
mem[16'hD116] = 8'hBD;
mem[16'hD117] = 8'h48;
mem[16'hD118] = 8'h50;
mem[16'hD119] = 8'h4C;
mem[16'hD11A] = 8'h4F;
mem[16'hD11B] = 8'hD4;
mem[16'hD11C] = 8'h44;
mem[16'hD11D] = 8'h52;
mem[16'hD11E] = 8'h41;
mem[16'hD11F] = 8'hD7;
mem[16'hD120] = 8'h58;
mem[16'hD121] = 8'h44;
mem[16'hD122] = 8'h52;
mem[16'hD123] = 8'h41;
mem[16'hD124] = 8'hD7;
mem[16'hD125] = 8'h48;
mem[16'hD126] = 8'h54;
mem[16'hD127] = 8'h41;
mem[16'hD128] = 8'hC2;
mem[16'hD129] = 8'h48;
mem[16'hD12A] = 8'h4F;
mem[16'hD12B] = 8'h4D;
mem[16'hD12C] = 8'hC5;
mem[16'hD12D] = 8'h52;
mem[16'hD12E] = 8'h4F;
mem[16'hD12F] = 8'h54;
mem[16'hD130] = 8'hBD;
mem[16'hD131] = 8'h53;
mem[16'hD132] = 8'h43;
mem[16'hD133] = 8'h41;
mem[16'hD134] = 8'h4C;
mem[16'hD135] = 8'h45;
mem[16'hD136] = 8'hBD;
mem[16'hD137] = 8'h53;
mem[16'hD138] = 8'h48;
mem[16'hD139] = 8'h4C;
mem[16'hD13A] = 8'h4F;
mem[16'hD13B] = 8'h41;
mem[16'hD13C] = 8'hC4;
mem[16'hD13D] = 8'h54;
mem[16'hD13E] = 8'h52;
mem[16'hD13F] = 8'h41;
mem[16'hD140] = 8'h43;
mem[16'hD141] = 8'hC5;
mem[16'hD142] = 8'h4E;
mem[16'hD143] = 8'h4F;
mem[16'hD144] = 8'h54;
mem[16'hD145] = 8'h52;
mem[16'hD146] = 8'h41;
mem[16'hD147] = 8'h43;
mem[16'hD148] = 8'hC5;
mem[16'hD149] = 8'h4E;
mem[16'hD14A] = 8'h4F;
mem[16'hD14B] = 8'h52;
mem[16'hD14C] = 8'h4D;
mem[16'hD14D] = 8'h41;
mem[16'hD14E] = 8'hCC;
mem[16'hD14F] = 8'h49;
mem[16'hD150] = 8'h4E;
mem[16'hD151] = 8'h56;
mem[16'hD152] = 8'h45;
mem[16'hD153] = 8'h52;
mem[16'hD154] = 8'h53;
mem[16'hD155] = 8'hC5;
mem[16'hD156] = 8'h46;
mem[16'hD157] = 8'h4C;
mem[16'hD158] = 8'h41;
mem[16'hD159] = 8'h53;
mem[16'hD15A] = 8'hC8;
mem[16'hD15B] = 8'h43;
mem[16'hD15C] = 8'h4F;
mem[16'hD15D] = 8'h4C;
mem[16'hD15E] = 8'h4F;
mem[16'hD15F] = 8'h52;
mem[16'hD160] = 8'hBD;
mem[16'hD161] = 8'h50;
mem[16'hD162] = 8'h4F;
mem[16'hD163] = 8'hD0;
mem[16'hD164] = 8'h56;
mem[16'hD165] = 8'h54;
mem[16'hD166] = 8'h41;
mem[16'hD167] = 8'hC2;
mem[16'hD168] = 8'h48;
mem[16'hD169] = 8'h49;
mem[16'hD16A] = 8'h4D;
mem[16'hD16B] = 8'h45;
mem[16'hD16C] = 8'h4D;
mem[16'hD16D] = 8'hBA;
mem[16'hD16E] = 8'h4C;
mem[16'hD16F] = 8'h4F;
mem[16'hD170] = 8'h4D;
mem[16'hD171] = 8'h45;
mem[16'hD172] = 8'h4D;
mem[16'hD173] = 8'hBA;
mem[16'hD174] = 8'h4F;
mem[16'hD175] = 8'h4E;
mem[16'hD176] = 8'h45;
mem[16'hD177] = 8'h52;
mem[16'hD178] = 8'hD2;
mem[16'hD179] = 8'h52;
mem[16'hD17A] = 8'h45;
mem[16'hD17B] = 8'h53;
mem[16'hD17C] = 8'h55;
mem[16'hD17D] = 8'h4D;
mem[16'hD17E] = 8'hC5;
mem[16'hD17F] = 8'h52;
mem[16'hD180] = 8'h45;
mem[16'hD181] = 8'h43;
mem[16'hD182] = 8'h41;
mem[16'hD183] = 8'h4C;
mem[16'hD184] = 8'hCC;
mem[16'hD185] = 8'h53;
mem[16'hD186] = 8'h54;
mem[16'hD187] = 8'h4F;
mem[16'hD188] = 8'h52;
mem[16'hD189] = 8'hC5;
mem[16'hD18A] = 8'h53;
mem[16'hD18B] = 8'h50;
mem[16'hD18C] = 8'h45;
mem[16'hD18D] = 8'h45;
mem[16'hD18E] = 8'h44;
mem[16'hD18F] = 8'hBD;
mem[16'hD190] = 8'h4C;
mem[16'hD191] = 8'h45;
mem[16'hD192] = 8'hD4;
mem[16'hD193] = 8'h47;
mem[16'hD194] = 8'h4F;
mem[16'hD195] = 8'h54;
mem[16'hD196] = 8'hCF;
mem[16'hD197] = 8'h52;
mem[16'hD198] = 8'h55;
mem[16'hD199] = 8'hCE;
mem[16'hD19A] = 8'h49;
mem[16'hD19B] = 8'hC6;
mem[16'hD19C] = 8'h52;
mem[16'hD19D] = 8'h45;
mem[16'hD19E] = 8'h53;
mem[16'hD19F] = 8'h54;
mem[16'hD1A0] = 8'h4F;
mem[16'hD1A1] = 8'h52;
mem[16'hD1A2] = 8'hC5;
mem[16'hD1A3] = 8'hA6;
mem[16'hD1A4] = 8'h47;
mem[16'hD1A5] = 8'h4F;
mem[16'hD1A6] = 8'h53;
mem[16'hD1A7] = 8'h55;
mem[16'hD1A8] = 8'hC2;
mem[16'hD1A9] = 8'h52;
mem[16'hD1AA] = 8'h45;
mem[16'hD1AB] = 8'h54;
mem[16'hD1AC] = 8'h55;
mem[16'hD1AD] = 8'h52;
mem[16'hD1AE] = 8'hCE;
mem[16'hD1AF] = 8'h52;
mem[16'hD1B0] = 8'h45;
mem[16'hD1B1] = 8'hCD;
mem[16'hD1B2] = 8'h53;
mem[16'hD1B3] = 8'h54;
mem[16'hD1B4] = 8'h4F;
mem[16'hD1B5] = 8'hD0;
mem[16'hD1B6] = 8'h4F;
mem[16'hD1B7] = 8'hCE;
mem[16'hD1B8] = 8'h57;
mem[16'hD1B9] = 8'h41;
mem[16'hD1BA] = 8'h49;
mem[16'hD1BB] = 8'hD4;
mem[16'hD1BC] = 8'h4C;
mem[16'hD1BD] = 8'h4F;
mem[16'hD1BE] = 8'h41;
mem[16'hD1BF] = 8'hC4;
mem[16'hD1C0] = 8'h53;
mem[16'hD1C1] = 8'h41;
mem[16'hD1C2] = 8'h56;
mem[16'hD1C3] = 8'hC5;
mem[16'hD1C4] = 8'h44;
mem[16'hD1C5] = 8'h45;
mem[16'hD1C6] = 8'hC6;
mem[16'hD1C7] = 8'h50;
mem[16'hD1C8] = 8'h4F;
mem[16'hD1C9] = 8'h4B;
mem[16'hD1CA] = 8'hC5;
mem[16'hD1CB] = 8'h50;
mem[16'hD1CC] = 8'h52;
mem[16'hD1CD] = 8'h49;
mem[16'hD1CE] = 8'h4E;
mem[16'hD1CF] = 8'hD4;
mem[16'hD1D0] = 8'h43;
mem[16'hD1D1] = 8'h4F;
mem[16'hD1D2] = 8'h4E;
mem[16'hD1D3] = 8'hD4;
mem[16'hD1D4] = 8'h4C;
mem[16'hD1D5] = 8'h49;
mem[16'hD1D6] = 8'h53;
mem[16'hD1D7] = 8'hD4;
mem[16'hD1D8] = 8'h43;
mem[16'hD1D9] = 8'h4C;
mem[16'hD1DA] = 8'h45;
mem[16'hD1DB] = 8'h41;
mem[16'hD1DC] = 8'hD2;
mem[16'hD1DD] = 8'h47;
mem[16'hD1DE] = 8'h45;
mem[16'hD1DF] = 8'hD4;
mem[16'hD1E0] = 8'h4E;
mem[16'hD1E1] = 8'h45;
mem[16'hD1E2] = 8'hD7;
mem[16'hD1E3] = 8'h54;
mem[16'hD1E4] = 8'h41;
mem[16'hD1E5] = 8'h42;
mem[16'hD1E6] = 8'hA8;
mem[16'hD1E7] = 8'h54;
mem[16'hD1E8] = 8'hCF;
mem[16'hD1E9] = 8'h46;
mem[16'hD1EA] = 8'hCE;
mem[16'hD1EB] = 8'h53;
mem[16'hD1EC] = 8'h50;
mem[16'hD1ED] = 8'h43;
mem[16'hD1EE] = 8'hA8;
mem[16'hD1EF] = 8'h54;
mem[16'hD1F0] = 8'h48;
mem[16'hD1F1] = 8'h45;
mem[16'hD1F2] = 8'hCE;
mem[16'hD1F3] = 8'h41;
mem[16'hD1F4] = 8'hD4;
mem[16'hD1F5] = 8'h4E;
mem[16'hD1F6] = 8'h4F;
mem[16'hD1F7] = 8'hD4;
mem[16'hD1F8] = 8'h53;
mem[16'hD1F9] = 8'h54;
mem[16'hD1FA] = 8'h45;
mem[16'hD1FB] = 8'hD0;
mem[16'hD1FC] = 8'hAB;
mem[16'hD1FD] = 8'hAD;
mem[16'hD1FE] = 8'hAA;
mem[16'hD1FF] = 8'hAF;
mem[16'hD200] = 8'hDE;
mem[16'hD201] = 8'h41;
mem[16'hD202] = 8'h4E;
mem[16'hD203] = 8'hC4;
mem[16'hD204] = 8'h4F;
mem[16'hD205] = 8'hD2;
mem[16'hD206] = 8'hBE;
mem[16'hD207] = 8'hBD;
mem[16'hD208] = 8'hBC;
mem[16'hD209] = 8'h53;
mem[16'hD20A] = 8'h47;
mem[16'hD20B] = 8'hCE;
mem[16'hD20C] = 8'h49;
mem[16'hD20D] = 8'h4E;
mem[16'hD20E] = 8'hD4;
mem[16'hD20F] = 8'h41;
mem[16'hD210] = 8'h42;
mem[16'hD211] = 8'hD3;
mem[16'hD212] = 8'h55;
mem[16'hD213] = 8'h53;
mem[16'hD214] = 8'hD2;
mem[16'hD215] = 8'h46;
mem[16'hD216] = 8'h52;
mem[16'hD217] = 8'hC5;
mem[16'hD218] = 8'h53;
mem[16'hD219] = 8'h43;
mem[16'hD21A] = 8'h52;
mem[16'hD21B] = 8'h4E;
mem[16'hD21C] = 8'hA8;
mem[16'hD21D] = 8'h50;
mem[16'hD21E] = 8'h44;
mem[16'hD21F] = 8'hCC;
mem[16'hD220] = 8'h50;
mem[16'hD221] = 8'h4F;
mem[16'hD222] = 8'hD3;
mem[16'hD223] = 8'h53;
mem[16'hD224] = 8'h51;
mem[16'hD225] = 8'hD2;
mem[16'hD226] = 8'h52;
mem[16'hD227] = 8'h4E;
mem[16'hD228] = 8'hC4;
mem[16'hD229] = 8'h4C;
mem[16'hD22A] = 8'h4F;
mem[16'hD22B] = 8'hC7;
mem[16'hD22C] = 8'h45;
mem[16'hD22D] = 8'h58;
mem[16'hD22E] = 8'hD0;
mem[16'hD22F] = 8'h43;
mem[16'hD230] = 8'h4F;
mem[16'hD231] = 8'hD3;
mem[16'hD232] = 8'h53;
mem[16'hD233] = 8'h49;
mem[16'hD234] = 8'hCE;
mem[16'hD235] = 8'h54;
mem[16'hD236] = 8'h41;
mem[16'hD237] = 8'hCE;
mem[16'hD238] = 8'h41;
mem[16'hD239] = 8'h54;
mem[16'hD23A] = 8'hCE;
mem[16'hD23B] = 8'h50;
mem[16'hD23C] = 8'h45;
mem[16'hD23D] = 8'h45;
mem[16'hD23E] = 8'hCB;
mem[16'hD23F] = 8'h4C;
mem[16'hD240] = 8'h45;
mem[16'hD241] = 8'hCE;
mem[16'hD242] = 8'h53;
mem[16'hD243] = 8'h54;
mem[16'hD244] = 8'h52;
mem[16'hD245] = 8'hA4;
mem[16'hD246] = 8'h56;
mem[16'hD247] = 8'h41;
mem[16'hD248] = 8'hCC;
mem[16'hD249] = 8'h41;
mem[16'hD24A] = 8'h53;
mem[16'hD24B] = 8'hC3;
mem[16'hD24C] = 8'h43;
mem[16'hD24D] = 8'h48;
mem[16'hD24E] = 8'h52;
mem[16'hD24F] = 8'hA4;
mem[16'hD250] = 8'h4C;
mem[16'hD251] = 8'h45;
mem[16'hD252] = 8'h46;
mem[16'hD253] = 8'h54;
mem[16'hD254] = 8'hA4;
mem[16'hD255] = 8'h52;
mem[16'hD256] = 8'h49;
mem[16'hD257] = 8'h47;
mem[16'hD258] = 8'h48;
mem[16'hD259] = 8'h54;
mem[16'hD25A] = 8'hA4;
mem[16'hD25B] = 8'h4D;
mem[16'hD25C] = 8'h49;
mem[16'hD25D] = 8'h44;
mem[16'hD25E] = 8'hA4;
mem[16'hD25F] = 8'h00;
mem[16'hD260] = 8'h4E;
mem[16'hD261] = 8'h45;
mem[16'hD262] = 8'h58;
mem[16'hD263] = 8'h54;
mem[16'hD264] = 8'h20;
mem[16'hD265] = 8'h57;
mem[16'hD266] = 8'h49;
mem[16'hD267] = 8'h54;
mem[16'hD268] = 8'h48;
mem[16'hD269] = 8'h4F;
mem[16'hD26A] = 8'h55;
mem[16'hD26B] = 8'h54;
mem[16'hD26C] = 8'h20;
mem[16'hD26D] = 8'h46;
mem[16'hD26E] = 8'h4F;
mem[16'hD26F] = 8'hD2;
mem[16'hD270] = 8'h53;
mem[16'hD271] = 8'h59;
mem[16'hD272] = 8'h4E;
mem[16'hD273] = 8'h54;
mem[16'hD274] = 8'h41;
mem[16'hD275] = 8'hD8;
mem[16'hD276] = 8'h52;
mem[16'hD277] = 8'h45;
mem[16'hD278] = 8'h54;
mem[16'hD279] = 8'h55;
mem[16'hD27A] = 8'h52;
mem[16'hD27B] = 8'h4E;
mem[16'hD27C] = 8'h20;
mem[16'hD27D] = 8'h57;
mem[16'hD27E] = 8'h49;
mem[16'hD27F] = 8'h54;
mem[16'hD280] = 8'h48;
mem[16'hD281] = 8'h4F;
mem[16'hD282] = 8'h55;
mem[16'hD283] = 8'h54;
mem[16'hD284] = 8'h20;
mem[16'hD285] = 8'h47;
mem[16'hD286] = 8'h4F;
mem[16'hD287] = 8'h53;
mem[16'hD288] = 8'h55;
mem[16'hD289] = 8'hC2;
mem[16'hD28A] = 8'h4F;
mem[16'hD28B] = 8'h55;
mem[16'hD28C] = 8'h54;
mem[16'hD28D] = 8'h20;
mem[16'hD28E] = 8'h4F;
mem[16'hD28F] = 8'h46;
mem[16'hD290] = 8'h20;
mem[16'hD291] = 8'h44;
mem[16'hD292] = 8'h41;
mem[16'hD293] = 8'h54;
mem[16'hD294] = 8'hC1;
mem[16'hD295] = 8'h49;
mem[16'hD296] = 8'h4C;
mem[16'hD297] = 8'h4C;
mem[16'hD298] = 8'h45;
mem[16'hD299] = 8'h47;
mem[16'hD29A] = 8'h41;
mem[16'hD29B] = 8'h4C;
mem[16'hD29C] = 8'h20;
mem[16'hD29D] = 8'h51;
mem[16'hD29E] = 8'h55;
mem[16'hD29F] = 8'h41;
mem[16'hD2A0] = 8'h4E;
mem[16'hD2A1] = 8'h54;
mem[16'hD2A2] = 8'h49;
mem[16'hD2A3] = 8'h54;
mem[16'hD2A4] = 8'hD9;
mem[16'hD2A5] = 8'h4F;
mem[16'hD2A6] = 8'h56;
mem[16'hD2A7] = 8'h45;
mem[16'hD2A8] = 8'h52;
mem[16'hD2A9] = 8'h46;
mem[16'hD2AA] = 8'h4C;
mem[16'hD2AB] = 8'h4F;
mem[16'hD2AC] = 8'hD7;
mem[16'hD2AD] = 8'h4F;
mem[16'hD2AE] = 8'h55;
mem[16'hD2AF] = 8'h54;
mem[16'hD2B0] = 8'h20;
mem[16'hD2B1] = 8'h4F;
mem[16'hD2B2] = 8'h46;
mem[16'hD2B3] = 8'h20;
mem[16'hD2B4] = 8'h4D;
mem[16'hD2B5] = 8'h45;
mem[16'hD2B6] = 8'h4D;
mem[16'hD2B7] = 8'h4F;
mem[16'hD2B8] = 8'h52;
mem[16'hD2B9] = 8'hD9;
mem[16'hD2BA] = 8'h55;
mem[16'hD2BB] = 8'h4E;
mem[16'hD2BC] = 8'h44;
mem[16'hD2BD] = 8'h45;
mem[16'hD2BE] = 8'h46;
mem[16'hD2BF] = 8'h27;
mem[16'hD2C0] = 8'h44;
mem[16'hD2C1] = 8'h20;
mem[16'hD2C2] = 8'h53;
mem[16'hD2C3] = 8'h54;
mem[16'hD2C4] = 8'h41;
mem[16'hD2C5] = 8'h54;
mem[16'hD2C6] = 8'h45;
mem[16'hD2C7] = 8'h4D;
mem[16'hD2C8] = 8'h45;
mem[16'hD2C9] = 8'h4E;
mem[16'hD2CA] = 8'hD4;
mem[16'hD2CB] = 8'h42;
mem[16'hD2CC] = 8'h41;
mem[16'hD2CD] = 8'h44;
mem[16'hD2CE] = 8'h20;
mem[16'hD2CF] = 8'h53;
mem[16'hD2D0] = 8'h55;
mem[16'hD2D1] = 8'h42;
mem[16'hD2D2] = 8'h53;
mem[16'hD2D3] = 8'h43;
mem[16'hD2D4] = 8'h52;
mem[16'hD2D5] = 8'h49;
mem[16'hD2D6] = 8'h50;
mem[16'hD2D7] = 8'hD4;
mem[16'hD2D8] = 8'h52;
mem[16'hD2D9] = 8'h45;
mem[16'hD2DA] = 8'h44;
mem[16'hD2DB] = 8'h49;
mem[16'hD2DC] = 8'h4D;
mem[16'hD2DD] = 8'h27;
mem[16'hD2DE] = 8'h44;
mem[16'hD2DF] = 8'h20;
mem[16'hD2E0] = 8'h41;
mem[16'hD2E1] = 8'h52;
mem[16'hD2E2] = 8'h52;
mem[16'hD2E3] = 8'h41;
mem[16'hD2E4] = 8'hD9;
mem[16'hD2E5] = 8'h44;
mem[16'hD2E6] = 8'h49;
mem[16'hD2E7] = 8'h56;
mem[16'hD2E8] = 8'h49;
mem[16'hD2E9] = 8'h53;
mem[16'hD2EA] = 8'h49;
mem[16'hD2EB] = 8'h4F;
mem[16'hD2EC] = 8'h4E;
mem[16'hD2ED] = 8'h20;
mem[16'hD2EE] = 8'h42;
mem[16'hD2EF] = 8'h59;
mem[16'hD2F0] = 8'h20;
mem[16'hD2F1] = 8'h5A;
mem[16'hD2F2] = 8'h45;
mem[16'hD2F3] = 8'h52;
mem[16'hD2F4] = 8'hCF;
mem[16'hD2F5] = 8'h49;
mem[16'hD2F6] = 8'h4C;
mem[16'hD2F7] = 8'h4C;
mem[16'hD2F8] = 8'h45;
mem[16'hD2F9] = 8'h47;
mem[16'hD2FA] = 8'h41;
mem[16'hD2FB] = 8'h4C;
mem[16'hD2FC] = 8'h20;
mem[16'hD2FD] = 8'h44;
mem[16'hD2FE] = 8'h49;
mem[16'hD2FF] = 8'h52;
mem[16'hD300] = 8'h45;
mem[16'hD301] = 8'h43;
mem[16'hD302] = 8'hD4;
mem[16'hD303] = 8'h54;
mem[16'hD304] = 8'h59;
mem[16'hD305] = 8'h50;
mem[16'hD306] = 8'h45;
mem[16'hD307] = 8'h20;
mem[16'hD308] = 8'h4D;
mem[16'hD309] = 8'h49;
mem[16'hD30A] = 8'h53;
mem[16'hD30B] = 8'h4D;
mem[16'hD30C] = 8'h41;
mem[16'hD30D] = 8'h54;
mem[16'hD30E] = 8'h43;
mem[16'hD30F] = 8'hC8;
mem[16'hD310] = 8'h53;
mem[16'hD311] = 8'h54;
mem[16'hD312] = 8'h52;
mem[16'hD313] = 8'h49;
mem[16'hD314] = 8'h4E;
mem[16'hD315] = 8'h47;
mem[16'hD316] = 8'h20;
mem[16'hD317] = 8'h54;
mem[16'hD318] = 8'h4F;
mem[16'hD319] = 8'h4F;
mem[16'hD31A] = 8'h20;
mem[16'hD31B] = 8'h4C;
mem[16'hD31C] = 8'h4F;
mem[16'hD31D] = 8'h4E;
mem[16'hD31E] = 8'hC7;
mem[16'hD31F] = 8'h46;
mem[16'hD320] = 8'h4F;
mem[16'hD321] = 8'h52;
mem[16'hD322] = 8'h4D;
mem[16'hD323] = 8'h55;
mem[16'hD324] = 8'h4C;
mem[16'hD325] = 8'h41;
mem[16'hD326] = 8'h20;
mem[16'hD327] = 8'h54;
mem[16'hD328] = 8'h4F;
mem[16'hD329] = 8'h4F;
mem[16'hD32A] = 8'h20;
mem[16'hD32B] = 8'h43;
mem[16'hD32C] = 8'h4F;
mem[16'hD32D] = 8'h4D;
mem[16'hD32E] = 8'h50;
mem[16'hD32F] = 8'h4C;
mem[16'hD330] = 8'h45;
mem[16'hD331] = 8'hD8;
mem[16'hD332] = 8'h43;
mem[16'hD333] = 8'h41;
mem[16'hD334] = 8'h4E;
mem[16'hD335] = 8'h27;
mem[16'hD336] = 8'h54;
mem[16'hD337] = 8'h20;
mem[16'hD338] = 8'h43;
mem[16'hD339] = 8'h4F;
mem[16'hD33A] = 8'h4E;
mem[16'hD33B] = 8'h54;
mem[16'hD33C] = 8'h49;
mem[16'hD33D] = 8'h4E;
mem[16'hD33E] = 8'h55;
mem[16'hD33F] = 8'hC5;
mem[16'hD340] = 8'h55;
mem[16'hD341] = 8'h4E;
mem[16'hD342] = 8'h44;
mem[16'hD343] = 8'h45;
mem[16'hD344] = 8'h46;
mem[16'hD345] = 8'h27;
mem[16'hD346] = 8'h44;
mem[16'hD347] = 8'h20;
mem[16'hD348] = 8'h46;
mem[16'hD349] = 8'h55;
mem[16'hD34A] = 8'h4E;
mem[16'hD34B] = 8'h43;
mem[16'hD34C] = 8'h54;
mem[16'hD34D] = 8'h49;
mem[16'hD34E] = 8'h4F;
mem[16'hD34F] = 8'hCE;
mem[16'hD350] = 8'h20;
mem[16'hD351] = 8'h45;
mem[16'hD352] = 8'h52;
mem[16'hD353] = 8'h52;
mem[16'hD354] = 8'h4F;
mem[16'hD355] = 8'h52;
mem[16'hD356] = 8'h07;
mem[16'hD357] = 8'h00;
mem[16'hD358] = 8'h20;
mem[16'hD359] = 8'h49;
mem[16'hD35A] = 8'h4E;
mem[16'hD35B] = 8'h20;
mem[16'hD35C] = 8'h00;
mem[16'hD35D] = 8'h0D;
mem[16'hD35E] = 8'h42;
mem[16'hD35F] = 8'h52;
mem[16'hD360] = 8'h45;
mem[16'hD361] = 8'h41;
mem[16'hD362] = 8'h4B;
mem[16'hD363] = 8'h07;
mem[16'hD364] = 8'h00;
mem[16'hD365] = 8'hBA;
mem[16'hD366] = 8'hE8;
mem[16'hD367] = 8'hE8;
mem[16'hD368] = 8'hE8;
mem[16'hD369] = 8'hE8;
mem[16'hD36A] = 8'hBD;
mem[16'hD36B] = 8'h01;
mem[16'hD36C] = 8'h01;
mem[16'hD36D] = 8'hC9;
mem[16'hD36E] = 8'h81;
mem[16'hD36F] = 8'hD0;
mem[16'hD370] = 8'h21;
mem[16'hD371] = 8'hA5;
mem[16'hD372] = 8'h86;
mem[16'hD373] = 8'hD0;
mem[16'hD374] = 8'h0A;
mem[16'hD375] = 8'hBD;
mem[16'hD376] = 8'h02;
mem[16'hD377] = 8'h01;
mem[16'hD378] = 8'h85;
mem[16'hD379] = 8'h85;
mem[16'hD37A] = 8'hBD;
mem[16'hD37B] = 8'h03;
mem[16'hD37C] = 8'h01;
mem[16'hD37D] = 8'h85;
mem[16'hD37E] = 8'h86;
mem[16'hD37F] = 8'hDD;
mem[16'hD380] = 8'h03;
mem[16'hD381] = 8'h01;
mem[16'hD382] = 8'hD0;
mem[16'hD383] = 8'h07;
mem[16'hD384] = 8'hA5;
mem[16'hD385] = 8'h85;
mem[16'hD386] = 8'hDD;
mem[16'hD387] = 8'h02;
mem[16'hD388] = 8'h01;
mem[16'hD389] = 8'hF0;
mem[16'hD38A] = 8'h07;
mem[16'hD38B] = 8'h8A;
mem[16'hD38C] = 8'h18;
mem[16'hD38D] = 8'h69;
mem[16'hD38E] = 8'h12;
mem[16'hD38F] = 8'hAA;
mem[16'hD390] = 8'hD0;
mem[16'hD391] = 8'hD8;
mem[16'hD392] = 8'h60;
mem[16'hD393] = 8'h20;
mem[16'hD394] = 8'hE3;
mem[16'hD395] = 8'hD3;
mem[16'hD396] = 8'h85;
mem[16'hD397] = 8'h6D;
mem[16'hD398] = 8'h84;
mem[16'hD399] = 8'h6E;
mem[16'hD39A] = 8'h38;
mem[16'hD39B] = 8'hA5;
mem[16'hD39C] = 8'h96;
mem[16'hD39D] = 8'hE5;
mem[16'hD39E] = 8'h9B;
mem[16'hD39F] = 8'h85;
mem[16'hD3A0] = 8'h5E;
mem[16'hD3A1] = 8'hA8;
mem[16'hD3A2] = 8'hA5;
mem[16'hD3A3] = 8'h97;
mem[16'hD3A4] = 8'hE5;
mem[16'hD3A5] = 8'h9C;
mem[16'hD3A6] = 8'hAA;
mem[16'hD3A7] = 8'hE8;
mem[16'hD3A8] = 8'h98;
mem[16'hD3A9] = 8'hF0;
mem[16'hD3AA] = 8'h23;
mem[16'hD3AB] = 8'hA5;
mem[16'hD3AC] = 8'h96;
mem[16'hD3AD] = 8'h38;
mem[16'hD3AE] = 8'hE5;
mem[16'hD3AF] = 8'h5E;
mem[16'hD3B0] = 8'h85;
mem[16'hD3B1] = 8'h96;
mem[16'hD3B2] = 8'hB0;
mem[16'hD3B3] = 8'h03;
mem[16'hD3B4] = 8'hC6;
mem[16'hD3B5] = 8'h97;
mem[16'hD3B6] = 8'h38;
mem[16'hD3B7] = 8'hA5;
mem[16'hD3B8] = 8'h94;
mem[16'hD3B9] = 8'hE5;
mem[16'hD3BA] = 8'h5E;
mem[16'hD3BB] = 8'h85;
mem[16'hD3BC] = 8'h94;
mem[16'hD3BD] = 8'hB0;
mem[16'hD3BE] = 8'h08;
mem[16'hD3BF] = 8'hC6;
mem[16'hD3C0] = 8'h95;
mem[16'hD3C1] = 8'h90;
mem[16'hD3C2] = 8'h04;
mem[16'hD3C3] = 8'hB1;
mem[16'hD3C4] = 8'h96;
mem[16'hD3C5] = 8'h91;
mem[16'hD3C6] = 8'h94;
mem[16'hD3C7] = 8'h88;
mem[16'hD3C8] = 8'hD0;
mem[16'hD3C9] = 8'hF9;
mem[16'hD3CA] = 8'hB1;
mem[16'hD3CB] = 8'h96;
mem[16'hD3CC] = 8'h91;
mem[16'hD3CD] = 8'h94;
mem[16'hD3CE] = 8'hC6;
mem[16'hD3CF] = 8'h97;
mem[16'hD3D0] = 8'hC6;
mem[16'hD3D1] = 8'h95;
mem[16'hD3D2] = 8'hCA;
mem[16'hD3D3] = 8'hD0;
mem[16'hD3D4] = 8'hF2;
mem[16'hD3D5] = 8'h60;
mem[16'hD3D6] = 8'h0A;
mem[16'hD3D7] = 8'h69;
mem[16'hD3D8] = 8'h36;
mem[16'hD3D9] = 8'hB0;
mem[16'hD3DA] = 8'h35;
mem[16'hD3DB] = 8'h85;
mem[16'hD3DC] = 8'h5E;
mem[16'hD3DD] = 8'hBA;
mem[16'hD3DE] = 8'hE4;
mem[16'hD3DF] = 8'h5E;
mem[16'hD3E0] = 8'h90;
mem[16'hD3E1] = 8'h2E;
mem[16'hD3E2] = 8'h60;
mem[16'hD3E3] = 8'hC4;
mem[16'hD3E4] = 8'h70;
mem[16'hD3E5] = 8'h90;
mem[16'hD3E6] = 8'h28;
mem[16'hD3E7] = 8'hD0;
mem[16'hD3E8] = 8'h04;
mem[16'hD3E9] = 8'hC5;
mem[16'hD3EA] = 8'h6F;
mem[16'hD3EB] = 8'h90;
mem[16'hD3EC] = 8'h22;
mem[16'hD3ED] = 8'h48;
mem[16'hD3EE] = 8'hA2;
mem[16'hD3EF] = 8'h09;
mem[16'hD3F0] = 8'h98;
mem[16'hD3F1] = 8'h48;
mem[16'hD3F2] = 8'hB5;
mem[16'hD3F3] = 8'h93;
mem[16'hD3F4] = 8'hCA;
mem[16'hD3F5] = 8'h10;
mem[16'hD3F6] = 8'hFA;
mem[16'hD3F7] = 8'h20;
mem[16'hD3F8] = 8'h84;
mem[16'hD3F9] = 8'hE4;
mem[16'hD3FA] = 8'hA2;
mem[16'hD3FB] = 8'hF7;
mem[16'hD3FC] = 8'h68;
mem[16'hD3FD] = 8'h95;
mem[16'hD3FE] = 8'h9D;
mem[16'hD3FF] = 8'hE8;
mem[16'hD400] = 8'h30;
mem[16'hD401] = 8'hFA;
mem[16'hD402] = 8'h68;
mem[16'hD403] = 8'hA8;
mem[16'hD404] = 8'h68;
mem[16'hD405] = 8'hC4;
mem[16'hD406] = 8'h70;
mem[16'hD407] = 8'h90;
mem[16'hD408] = 8'h06;
mem[16'hD409] = 8'hD0;
mem[16'hD40A] = 8'h05;
mem[16'hD40B] = 8'hC5;
mem[16'hD40C] = 8'h6F;
mem[16'hD40D] = 8'hB0;
mem[16'hD40E] = 8'h01;
mem[16'hD40F] = 8'h60;
mem[16'hD410] = 8'hA2;
mem[16'hD411] = 8'h4D;
mem[16'hD412] = 8'h24;
mem[16'hD413] = 8'hD8;
mem[16'hD414] = 8'h10;
mem[16'hD415] = 8'h03;
mem[16'hD416] = 8'h4C;
mem[16'hD417] = 8'hE9;
mem[16'hD418] = 8'hF2;
mem[16'hD419] = 8'h20;
mem[16'hD41A] = 8'hFB;
mem[16'hD41B] = 8'hDA;
mem[16'hD41C] = 8'h20;
mem[16'hD41D] = 8'h5A;
mem[16'hD41E] = 8'hDB;
mem[16'hD41F] = 8'hBD;
mem[16'hD420] = 8'h60;
mem[16'hD421] = 8'hD2;
mem[16'hD422] = 8'h48;
mem[16'hD423] = 8'h20;
mem[16'hD424] = 8'h5C;
mem[16'hD425] = 8'hDB;
mem[16'hD426] = 8'hE8;
mem[16'hD427] = 8'h68;
mem[16'hD428] = 8'h10;
mem[16'hD429] = 8'hF5;
mem[16'hD42A] = 8'h20;
mem[16'hD42B] = 8'h83;
mem[16'hD42C] = 8'hD6;
mem[16'hD42D] = 8'hA9;
mem[16'hD42E] = 8'h50;
mem[16'hD42F] = 8'hA0;
mem[16'hD430] = 8'hD3;
mem[16'hD431] = 8'h20;
mem[16'hD432] = 8'h3A;
mem[16'hD433] = 8'hDB;
mem[16'hD434] = 8'hA4;
mem[16'hD435] = 8'h76;
mem[16'hD436] = 8'hC8;
mem[16'hD437] = 8'hF0;
mem[16'hD438] = 8'h03;
mem[16'hD439] = 8'h20;
mem[16'hD43A] = 8'h19;
mem[16'hD43B] = 8'hED;
mem[16'hD43C] = 8'h20;
mem[16'hD43D] = 8'hFB;
mem[16'hD43E] = 8'hDA;
mem[16'hD43F] = 8'hA2;
mem[16'hD440] = 8'hDD;
mem[16'hD441] = 8'h20;
mem[16'hD442] = 8'h2E;
mem[16'hD443] = 8'hD5;
mem[16'hD444] = 8'h86;
mem[16'hD445] = 8'hB8;
mem[16'hD446] = 8'h84;
mem[16'hD447] = 8'hB9;
mem[16'hD448] = 8'h46;
mem[16'hD449] = 8'hD8;
mem[16'hD44A] = 8'h20;
mem[16'hD44B] = 8'hB1;
mem[16'hD44C] = 8'h00;
mem[16'hD44D] = 8'hAA;
mem[16'hD44E] = 8'hF0;
mem[16'hD44F] = 8'hEC;
mem[16'hD450] = 8'hA2;
mem[16'hD451] = 8'hFF;
mem[16'hD452] = 8'h86;
mem[16'hD453] = 8'h76;
mem[16'hD454] = 8'h90;
mem[16'hD455] = 8'h06;
mem[16'hD456] = 8'h20;
mem[16'hD457] = 8'h59;
mem[16'hD458] = 8'hD5;
mem[16'hD459] = 8'h4C;
mem[16'hD45A] = 8'h05;
mem[16'hD45B] = 8'hD8;
mem[16'hD45C] = 8'hA6;
mem[16'hD45D] = 8'hAF;
mem[16'hD45E] = 8'h86;
mem[16'hD45F] = 8'h69;
mem[16'hD460] = 8'hA6;
mem[16'hD461] = 8'hB0;
mem[16'hD462] = 8'h86;
mem[16'hD463] = 8'h6A;
mem[16'hD464] = 8'h20;
mem[16'hD465] = 8'h0C;
mem[16'hD466] = 8'hDA;
mem[16'hD467] = 8'h20;
mem[16'hD468] = 8'h59;
mem[16'hD469] = 8'hD5;
mem[16'hD46A] = 8'h84;
mem[16'hD46B] = 8'h0F;
mem[16'hD46C] = 8'h20;
mem[16'hD46D] = 8'h1A;
mem[16'hD46E] = 8'hD6;
mem[16'hD46F] = 8'h90;
mem[16'hD470] = 8'h44;
mem[16'hD471] = 8'hA0;
mem[16'hD472] = 8'h01;
mem[16'hD473] = 8'hB1;
mem[16'hD474] = 8'h9B;
mem[16'hD475] = 8'h85;
mem[16'hD476] = 8'h5F;
mem[16'hD477] = 8'hA5;
mem[16'hD478] = 8'h69;
mem[16'hD479] = 8'h85;
mem[16'hD47A] = 8'h5E;
mem[16'hD47B] = 8'hA5;
mem[16'hD47C] = 8'h9C;
mem[16'hD47D] = 8'h85;
mem[16'hD47E] = 8'h61;
mem[16'hD47F] = 8'hA5;
mem[16'hD480] = 8'h9B;
mem[16'hD481] = 8'h88;
mem[16'hD482] = 8'hF1;
mem[16'hD483] = 8'h9B;
mem[16'hD484] = 8'h18;
mem[16'hD485] = 8'h65;
mem[16'hD486] = 8'h69;
mem[16'hD487] = 8'h85;
mem[16'hD488] = 8'h69;
mem[16'hD489] = 8'h85;
mem[16'hD48A] = 8'h60;
mem[16'hD48B] = 8'hA5;
mem[16'hD48C] = 8'h6A;
mem[16'hD48D] = 8'h69;
mem[16'hD48E] = 8'hFF;
mem[16'hD48F] = 8'h85;
mem[16'hD490] = 8'h6A;
mem[16'hD491] = 8'hE5;
mem[16'hD492] = 8'h9C;
mem[16'hD493] = 8'hAA;
mem[16'hD494] = 8'h38;
mem[16'hD495] = 8'hA5;
mem[16'hD496] = 8'h9B;
mem[16'hD497] = 8'hE5;
mem[16'hD498] = 8'h69;
mem[16'hD499] = 8'hA8;
mem[16'hD49A] = 8'hB0;
mem[16'hD49B] = 8'h03;
mem[16'hD49C] = 8'hE8;
mem[16'hD49D] = 8'hC6;
mem[16'hD49E] = 8'h61;
mem[16'hD49F] = 8'h18;
mem[16'hD4A0] = 8'h65;
mem[16'hD4A1] = 8'h5E;
mem[16'hD4A2] = 8'h90;
mem[16'hD4A3] = 8'h03;
mem[16'hD4A4] = 8'hC6;
mem[16'hD4A5] = 8'h5F;
mem[16'hD4A6] = 8'h18;
mem[16'hD4A7] = 8'hB1;
mem[16'hD4A8] = 8'h5E;
mem[16'hD4A9] = 8'h91;
mem[16'hD4AA] = 8'h60;
mem[16'hD4AB] = 8'hC8;
mem[16'hD4AC] = 8'hD0;
mem[16'hD4AD] = 8'hF9;
mem[16'hD4AE] = 8'hE6;
mem[16'hD4AF] = 8'h5F;
mem[16'hD4B0] = 8'hE6;
mem[16'hD4B1] = 8'h61;
mem[16'hD4B2] = 8'hCA;
mem[16'hD4B3] = 8'hD0;
mem[16'hD4B4] = 8'hF2;
mem[16'hD4B5] = 8'hAD;
mem[16'hD4B6] = 8'h00;
mem[16'hD4B7] = 8'h02;
mem[16'hD4B8] = 8'hF0;
mem[16'hD4B9] = 8'h38;
mem[16'hD4BA] = 8'hA5;
mem[16'hD4BB] = 8'h73;
mem[16'hD4BC] = 8'hA4;
mem[16'hD4BD] = 8'h74;
mem[16'hD4BE] = 8'h85;
mem[16'hD4BF] = 8'h6F;
mem[16'hD4C0] = 8'h84;
mem[16'hD4C1] = 8'h70;
mem[16'hD4C2] = 8'hA5;
mem[16'hD4C3] = 8'h69;
mem[16'hD4C4] = 8'h85;
mem[16'hD4C5] = 8'h96;
mem[16'hD4C6] = 8'h65;
mem[16'hD4C7] = 8'h0F;
mem[16'hD4C8] = 8'h85;
mem[16'hD4C9] = 8'h94;
mem[16'hD4CA] = 8'hA4;
mem[16'hD4CB] = 8'h6A;
mem[16'hD4CC] = 8'h84;
mem[16'hD4CD] = 8'h97;
mem[16'hD4CE] = 8'h90;
mem[16'hD4CF] = 8'h01;
mem[16'hD4D0] = 8'hC8;
mem[16'hD4D1] = 8'h84;
mem[16'hD4D2] = 8'h95;
mem[16'hD4D3] = 8'h20;
mem[16'hD4D4] = 8'h93;
mem[16'hD4D5] = 8'hD3;
mem[16'hD4D6] = 8'hA5;
mem[16'hD4D7] = 8'h50;
mem[16'hD4D8] = 8'hA4;
mem[16'hD4D9] = 8'h51;
mem[16'hD4DA] = 8'h8D;
mem[16'hD4DB] = 8'hFE;
mem[16'hD4DC] = 8'h01;
mem[16'hD4DD] = 8'h8C;
mem[16'hD4DE] = 8'hFF;
mem[16'hD4DF] = 8'h01;
mem[16'hD4E0] = 8'hA5;
mem[16'hD4E1] = 8'h6D;
mem[16'hD4E2] = 8'hA4;
mem[16'hD4E3] = 8'h6E;
mem[16'hD4E4] = 8'h85;
mem[16'hD4E5] = 8'h69;
mem[16'hD4E6] = 8'h84;
mem[16'hD4E7] = 8'h6A;
mem[16'hD4E8] = 8'hA4;
mem[16'hD4E9] = 8'h0F;
mem[16'hD4EA] = 8'hB9;
mem[16'hD4EB] = 8'hFB;
mem[16'hD4EC] = 8'h01;
mem[16'hD4ED] = 8'h88;
mem[16'hD4EE] = 8'h91;
mem[16'hD4EF] = 8'h9B;
mem[16'hD4F0] = 8'hD0;
mem[16'hD4F1] = 8'hF8;
mem[16'hD4F2] = 8'h20;
mem[16'hD4F3] = 8'h65;
mem[16'hD4F4] = 8'hD6;
mem[16'hD4F5] = 8'hA5;
mem[16'hD4F6] = 8'h67;
mem[16'hD4F7] = 8'hA4;
mem[16'hD4F8] = 8'h68;
mem[16'hD4F9] = 8'h85;
mem[16'hD4FA] = 8'h5E;
mem[16'hD4FB] = 8'h84;
mem[16'hD4FC] = 8'h5F;
mem[16'hD4FD] = 8'h18;
mem[16'hD4FE] = 8'hA0;
mem[16'hD4FF] = 8'h01;
mem[16'hD500] = 8'hB1;
mem[16'hD501] = 8'h5E;
mem[16'hD502] = 8'hD0;
mem[16'hD503] = 8'h0B;
mem[16'hD504] = 8'hA5;
mem[16'hD505] = 8'h69;
mem[16'hD506] = 8'h85;
mem[16'hD507] = 8'hAF;
mem[16'hD508] = 8'hA5;
mem[16'hD509] = 8'h6A;
mem[16'hD50A] = 8'h85;
mem[16'hD50B] = 8'hB0;
mem[16'hD50C] = 8'h4C;
mem[16'hD50D] = 8'h3C;
mem[16'hD50E] = 8'hD4;
mem[16'hD50F] = 8'hA0;
mem[16'hD510] = 8'h04;
mem[16'hD511] = 8'hC8;
mem[16'hD512] = 8'hB1;
mem[16'hD513] = 8'h5E;
mem[16'hD514] = 8'hD0;
mem[16'hD515] = 8'hFB;
mem[16'hD516] = 8'hC8;
mem[16'hD517] = 8'h98;
mem[16'hD518] = 8'h65;
mem[16'hD519] = 8'h5E;
mem[16'hD51A] = 8'hAA;
mem[16'hD51B] = 8'hA0;
mem[16'hD51C] = 8'h00;
mem[16'hD51D] = 8'h91;
mem[16'hD51E] = 8'h5E;
mem[16'hD51F] = 8'hA5;
mem[16'hD520] = 8'h5F;
mem[16'hD521] = 8'h69;
mem[16'hD522] = 8'h00;
mem[16'hD523] = 8'hC8;
mem[16'hD524] = 8'h91;
mem[16'hD525] = 8'h5E;
mem[16'hD526] = 8'h86;
mem[16'hD527] = 8'h5E;
mem[16'hD528] = 8'h85;
mem[16'hD529] = 8'h5F;
mem[16'hD52A] = 8'h90;
mem[16'hD52B] = 8'hD2;
mem[16'hD52C] = 8'hA2;
mem[16'hD52D] = 8'h80;
mem[16'hD52E] = 8'h86;
mem[16'hD52F] = 8'h33;
mem[16'hD530] = 8'h20;
mem[16'hD531] = 8'h6A;
mem[16'hD532] = 8'hFD;
mem[16'hD533] = 8'hE0;
mem[16'hD534] = 8'hEF;
mem[16'hD535] = 8'h90;
mem[16'hD536] = 8'h02;
mem[16'hD537] = 8'hA2;
mem[16'hD538] = 8'hEF;
mem[16'hD539] = 8'hA9;
mem[16'hD53A] = 8'h00;
mem[16'hD53B] = 8'h9D;
mem[16'hD53C] = 8'h00;
mem[16'hD53D] = 8'h02;
mem[16'hD53E] = 8'h8A;
mem[16'hD53F] = 8'hF0;
mem[16'hD540] = 8'h0B;
mem[16'hD541] = 8'hBD;
mem[16'hD542] = 8'hFF;
mem[16'hD543] = 8'h01;
mem[16'hD544] = 8'h29;
mem[16'hD545] = 8'h7F;
mem[16'hD546] = 8'h9D;
mem[16'hD547] = 8'hFF;
mem[16'hD548] = 8'h01;
mem[16'hD549] = 8'hCA;
mem[16'hD54A] = 8'hD0;
mem[16'hD54B] = 8'hF5;
mem[16'hD54C] = 8'hA9;
mem[16'hD54D] = 8'h00;
mem[16'hD54E] = 8'hA2;
mem[16'hD54F] = 8'hFF;
mem[16'hD550] = 8'hA0;
mem[16'hD551] = 8'h01;
mem[16'hD552] = 8'h60;
mem[16'hD553] = 8'h20;
mem[16'hD554] = 8'h0C;
mem[16'hD555] = 8'hFD;
mem[16'hD556] = 8'h29;
mem[16'hD557] = 8'h7F;
mem[16'hD558] = 8'h60;
mem[16'hD559] = 8'hA6;
mem[16'hD55A] = 8'hB8;
mem[16'hD55B] = 8'hCA;
mem[16'hD55C] = 8'hA0;
mem[16'hD55D] = 8'h04;
mem[16'hD55E] = 8'h84;
mem[16'hD55F] = 8'h13;
mem[16'hD560] = 8'h24;
mem[16'hD561] = 8'hD6;
mem[16'hD562] = 8'h10;
mem[16'hD563] = 8'h08;
mem[16'hD564] = 8'h68;
mem[16'hD565] = 8'h68;
mem[16'hD566] = 8'h20;
mem[16'hD567] = 8'h65;
mem[16'hD568] = 8'hD6;
mem[16'hD569] = 8'h4C;
mem[16'hD56A] = 8'hD2;
mem[16'hD56B] = 8'hD7;
mem[16'hD56C] = 8'hE8;
mem[16'hD56D] = 8'hBD;
mem[16'hD56E] = 8'h00;
mem[16'hD56F] = 8'h02;
mem[16'hD570] = 8'h24;
mem[16'hD571] = 8'h13;
mem[16'hD572] = 8'h70;
mem[16'hD573] = 8'h04;
mem[16'hD574] = 8'hC9;
mem[16'hD575] = 8'h20;
mem[16'hD576] = 8'hF0;
mem[16'hD577] = 8'hF4;
mem[16'hD578] = 8'h85;
mem[16'hD579] = 8'h0E;
mem[16'hD57A] = 8'hC9;
mem[16'hD57B] = 8'h22;
mem[16'hD57C] = 8'hF0;
mem[16'hD57D] = 8'h74;
mem[16'hD57E] = 8'h70;
mem[16'hD57F] = 8'h4D;
mem[16'hD580] = 8'hC9;
mem[16'hD581] = 8'h3F;
mem[16'hD582] = 8'hD0;
mem[16'hD583] = 8'h04;
mem[16'hD584] = 8'hA9;
mem[16'hD585] = 8'hBA;
mem[16'hD586] = 8'hD0;
mem[16'hD587] = 8'h45;
mem[16'hD588] = 8'hC9;
mem[16'hD589] = 8'h30;
mem[16'hD58A] = 8'h90;
mem[16'hD58B] = 8'h04;
mem[16'hD58C] = 8'hC9;
mem[16'hD58D] = 8'h3C;
mem[16'hD58E] = 8'h90;
mem[16'hD58F] = 8'h3D;
mem[16'hD590] = 8'h84;
mem[16'hD591] = 8'hAD;
mem[16'hD592] = 8'hA9;
mem[16'hD593] = 8'hD0;
mem[16'hD594] = 8'h85;
mem[16'hD595] = 8'h9D;
mem[16'hD596] = 8'hA9;
mem[16'hD597] = 8'hCF;
mem[16'hD598] = 8'h85;
mem[16'hD599] = 8'h9E;
mem[16'hD59A] = 8'hA0;
mem[16'hD59B] = 8'h00;
mem[16'hD59C] = 8'h84;
mem[16'hD59D] = 8'h0F;
mem[16'hD59E] = 8'h88;
mem[16'hD59F] = 8'h86;
mem[16'hD5A0] = 8'hB8;
mem[16'hD5A1] = 8'hCA;
mem[16'hD5A2] = 8'hC8;
mem[16'hD5A3] = 8'hD0;
mem[16'hD5A4] = 8'h02;
mem[16'hD5A5] = 8'hE6;
mem[16'hD5A6] = 8'h9E;
mem[16'hD5A7] = 8'hE8;
mem[16'hD5A8] = 8'hBD;
mem[16'hD5A9] = 8'h00;
mem[16'hD5AA] = 8'h02;
mem[16'hD5AB] = 8'hC9;
mem[16'hD5AC] = 8'h20;
mem[16'hD5AD] = 8'hF0;
mem[16'hD5AE] = 8'hF8;
mem[16'hD5AF] = 8'h38;
mem[16'hD5B0] = 8'hF1;
mem[16'hD5B1] = 8'h9D;
mem[16'hD5B2] = 8'hF0;
mem[16'hD5B3] = 8'hEE;
mem[16'hD5B4] = 8'hC9;
mem[16'hD5B5] = 8'h80;
mem[16'hD5B6] = 8'hD0;
mem[16'hD5B7] = 8'h41;
mem[16'hD5B8] = 8'h05;
mem[16'hD5B9] = 8'h0F;
mem[16'hD5BA] = 8'hC9;
mem[16'hD5BB] = 8'hC5;
mem[16'hD5BC] = 8'hD0;
mem[16'hD5BD] = 8'h0D;
mem[16'hD5BE] = 8'hBD;
mem[16'hD5BF] = 8'h01;
mem[16'hD5C0] = 8'h02;
mem[16'hD5C1] = 8'hC9;
mem[16'hD5C2] = 8'h4E;
mem[16'hD5C3] = 8'hF0;
mem[16'hD5C4] = 8'h34;
mem[16'hD5C5] = 8'hC9;
mem[16'hD5C6] = 8'h4F;
mem[16'hD5C7] = 8'hF0;
mem[16'hD5C8] = 8'h30;
mem[16'hD5C9] = 8'hA9;
mem[16'hD5CA] = 8'hC5;
mem[16'hD5CB] = 8'hA4;
mem[16'hD5CC] = 8'hAD;
mem[16'hD5CD] = 8'hE8;
mem[16'hD5CE] = 8'hC8;
mem[16'hD5CF] = 8'h99;
mem[16'hD5D0] = 8'hFB;
mem[16'hD5D1] = 8'h01;
mem[16'hD5D2] = 8'hB9;
mem[16'hD5D3] = 8'hFB;
mem[16'hD5D4] = 8'h01;
mem[16'hD5D5] = 8'hF0;
mem[16'hD5D6] = 8'h39;
mem[16'hD5D7] = 8'h38;
mem[16'hD5D8] = 8'hE9;
mem[16'hD5D9] = 8'h3A;
mem[16'hD5DA] = 8'hF0;
mem[16'hD5DB] = 8'h04;
mem[16'hD5DC] = 8'hC9;
mem[16'hD5DD] = 8'h49;
mem[16'hD5DE] = 8'hD0;
mem[16'hD5DF] = 8'h02;
mem[16'hD5E0] = 8'h85;
mem[16'hD5E1] = 8'h13;
mem[16'hD5E2] = 8'h38;
mem[16'hD5E3] = 8'hE9;
mem[16'hD5E4] = 8'h78;
mem[16'hD5E5] = 8'hD0;
mem[16'hD5E6] = 8'h86;
mem[16'hD5E7] = 8'h85;
mem[16'hD5E8] = 8'h0E;
mem[16'hD5E9] = 8'hBD;
mem[16'hD5EA] = 8'h00;
mem[16'hD5EB] = 8'h02;
mem[16'hD5EC] = 8'hF0;
mem[16'hD5ED] = 8'hDF;
mem[16'hD5EE] = 8'hC5;
mem[16'hD5EF] = 8'h0E;
mem[16'hD5F0] = 8'hF0;
mem[16'hD5F1] = 8'hDB;
mem[16'hD5F2] = 8'hC8;
mem[16'hD5F3] = 8'h99;
mem[16'hD5F4] = 8'hFB;
mem[16'hD5F5] = 8'h01;
mem[16'hD5F6] = 8'hE8;
mem[16'hD5F7] = 8'hD0;
mem[16'hD5F8] = 8'hF0;
mem[16'hD5F9] = 8'hA6;
mem[16'hD5FA] = 8'hB8;
mem[16'hD5FB] = 8'hE6;
mem[16'hD5FC] = 8'h0F;
mem[16'hD5FD] = 8'hB1;
mem[16'hD5FE] = 8'h9D;
mem[16'hD5FF] = 8'hC8;
mem[16'hD600] = 8'hD0;
mem[16'hD601] = 8'h02;
mem[16'hD602] = 8'hE6;
mem[16'hD603] = 8'h9E;
mem[16'hD604] = 8'h0A;
mem[16'hD605] = 8'h90;
mem[16'hD606] = 8'hF6;
mem[16'hD607] = 8'hB1;
mem[16'hD608] = 8'h9D;
mem[16'hD609] = 8'hD0;
mem[16'hD60A] = 8'h9D;
mem[16'hD60B] = 8'hBD;
mem[16'hD60C] = 8'h00;
mem[16'hD60D] = 8'h02;
mem[16'hD60E] = 8'h10;
mem[16'hD60F] = 8'hBB;
mem[16'hD610] = 8'h99;
mem[16'hD611] = 8'hFD;
mem[16'hD612] = 8'h01;
mem[16'hD613] = 8'hC6;
mem[16'hD614] = 8'hB9;
mem[16'hD615] = 8'hA9;
mem[16'hD616] = 8'hFF;
mem[16'hD617] = 8'h85;
mem[16'hD618] = 8'hB8;
mem[16'hD619] = 8'h60;
mem[16'hD61A] = 8'hA5;
mem[16'hD61B] = 8'h67;
mem[16'hD61C] = 8'hA6;
mem[16'hD61D] = 8'h68;
mem[16'hD61E] = 8'hA0;
mem[16'hD61F] = 8'h01;
mem[16'hD620] = 8'h85;
mem[16'hD621] = 8'h9B;
mem[16'hD622] = 8'h86;
mem[16'hD623] = 8'h9C;
mem[16'hD624] = 8'hB1;
mem[16'hD625] = 8'h9B;
mem[16'hD626] = 8'hF0;
mem[16'hD627] = 8'h1F;
mem[16'hD628] = 8'hC8;
mem[16'hD629] = 8'hC8;
mem[16'hD62A] = 8'hA5;
mem[16'hD62B] = 8'h51;
mem[16'hD62C] = 8'hD1;
mem[16'hD62D] = 8'h9B;
mem[16'hD62E] = 8'h90;
mem[16'hD62F] = 8'h18;
mem[16'hD630] = 8'hF0;
mem[16'hD631] = 8'h03;
mem[16'hD632] = 8'h88;
mem[16'hD633] = 8'hD0;
mem[16'hD634] = 8'h09;
mem[16'hD635] = 8'hA5;
mem[16'hD636] = 8'h50;
mem[16'hD637] = 8'h88;
mem[16'hD638] = 8'hD1;
mem[16'hD639] = 8'h9B;
mem[16'hD63A] = 8'h90;
mem[16'hD63B] = 8'h0C;
mem[16'hD63C] = 8'hF0;
mem[16'hD63D] = 8'h0A;
mem[16'hD63E] = 8'h88;
mem[16'hD63F] = 8'hB1;
mem[16'hD640] = 8'h9B;
mem[16'hD641] = 8'hAA;
mem[16'hD642] = 8'h88;
mem[16'hD643] = 8'hB1;
mem[16'hD644] = 8'h9B;
mem[16'hD645] = 8'hB0;
mem[16'hD646] = 8'hD7;
mem[16'hD647] = 8'h18;
mem[16'hD648] = 8'h60;
mem[16'hD649] = 8'hD0;
mem[16'hD64A] = 8'hFD;
mem[16'hD64B] = 8'hA9;
mem[16'hD64C] = 8'h00;
mem[16'hD64D] = 8'h85;
mem[16'hD64E] = 8'hD6;
mem[16'hD64F] = 8'hA8;
mem[16'hD650] = 8'h91;
mem[16'hD651] = 8'h67;
mem[16'hD652] = 8'hC8;
mem[16'hD653] = 8'h91;
mem[16'hD654] = 8'h67;
mem[16'hD655] = 8'hA5;
mem[16'hD656] = 8'h67;
mem[16'hD657] = 8'h69;
mem[16'hD658] = 8'h02;
mem[16'hD659] = 8'h85;
mem[16'hD65A] = 8'h69;
mem[16'hD65B] = 8'h85;
mem[16'hD65C] = 8'hAF;
mem[16'hD65D] = 8'hA5;
mem[16'hD65E] = 8'h68;
mem[16'hD65F] = 8'h69;
mem[16'hD660] = 8'h00;
mem[16'hD661] = 8'h85;
mem[16'hD662] = 8'h6A;
mem[16'hD663] = 8'h85;
mem[16'hD664] = 8'hB0;
mem[16'hD665] = 8'h20;
mem[16'hD666] = 8'h97;
mem[16'hD667] = 8'hD6;
mem[16'hD668] = 8'hA9;
mem[16'hD669] = 8'h00;
mem[16'hD66A] = 8'hD0;
mem[16'hD66B] = 8'h2A;
mem[16'hD66C] = 8'hA5;
mem[16'hD66D] = 8'h73;
mem[16'hD66E] = 8'hA4;
mem[16'hD66F] = 8'h74;
mem[16'hD670] = 8'h85;
mem[16'hD671] = 8'h6F;
mem[16'hD672] = 8'h84;
mem[16'hD673] = 8'h70;
mem[16'hD674] = 8'hA5;
mem[16'hD675] = 8'h69;
mem[16'hD676] = 8'hA4;
mem[16'hD677] = 8'h6A;
mem[16'hD678] = 8'h85;
mem[16'hD679] = 8'h6B;
mem[16'hD67A] = 8'h84;
mem[16'hD67B] = 8'h6C;
mem[16'hD67C] = 8'h85;
mem[16'hD67D] = 8'h6D;
mem[16'hD67E] = 8'h84;
mem[16'hD67F] = 8'h6E;
mem[16'hD680] = 8'h20;
mem[16'hD681] = 8'h49;
mem[16'hD682] = 8'hD8;
mem[16'hD683] = 8'hA2;
mem[16'hD684] = 8'h55;
mem[16'hD685] = 8'h86;
mem[16'hD686] = 8'h52;
mem[16'hD687] = 8'h68;
mem[16'hD688] = 8'hA8;
mem[16'hD689] = 8'h68;
mem[16'hD68A] = 8'hA2;
mem[16'hD68B] = 8'hF8;
mem[16'hD68C] = 8'h9A;
mem[16'hD68D] = 8'h48;
mem[16'hD68E] = 8'h98;
mem[16'hD68F] = 8'h48;
mem[16'hD690] = 8'hA9;
mem[16'hD691] = 8'h00;
mem[16'hD692] = 8'h85;
mem[16'hD693] = 8'h7A;
mem[16'hD694] = 8'h85;
mem[16'hD695] = 8'h14;
mem[16'hD696] = 8'h60;
mem[16'hD697] = 8'h18;
mem[16'hD698] = 8'hA5;
mem[16'hD699] = 8'h67;
mem[16'hD69A] = 8'h69;
mem[16'hD69B] = 8'hFF;
mem[16'hD69C] = 8'h85;
mem[16'hD69D] = 8'hB8;
mem[16'hD69E] = 8'hA5;
mem[16'hD69F] = 8'h68;
mem[16'hD6A0] = 8'h69;
mem[16'hD6A1] = 8'hFF;
mem[16'hD6A2] = 8'h85;
mem[16'hD6A3] = 8'hB9;
mem[16'hD6A4] = 8'h60;
mem[16'hD6A5] = 8'h90;
mem[16'hD6A6] = 8'h0A;
mem[16'hD6A7] = 8'hF0;
mem[16'hD6A8] = 8'h08;
mem[16'hD6A9] = 8'hC9;
mem[16'hD6AA] = 8'hC9;
mem[16'hD6AB] = 8'hF0;
mem[16'hD6AC] = 8'h04;
mem[16'hD6AD] = 8'hC9;
mem[16'hD6AE] = 8'h2C;
mem[16'hD6AF] = 8'hD0;
mem[16'hD6B0] = 8'hE5;
mem[16'hD6B1] = 8'h20;
mem[16'hD6B2] = 8'h0C;
mem[16'hD6B3] = 8'hDA;
mem[16'hD6B4] = 8'h20;
mem[16'hD6B5] = 8'h1A;
mem[16'hD6B6] = 8'hD6;
mem[16'hD6B7] = 8'h20;
mem[16'hD6B8] = 8'hB7;
mem[16'hD6B9] = 8'h00;
mem[16'hD6BA] = 8'hF0;
mem[16'hD6BB] = 8'h10;
mem[16'hD6BC] = 8'hC9;
mem[16'hD6BD] = 8'hC9;
mem[16'hD6BE] = 8'hF0;
mem[16'hD6BF] = 8'h04;
mem[16'hD6C0] = 8'hC9;
mem[16'hD6C1] = 8'h2C;
mem[16'hD6C2] = 8'hD0;
mem[16'hD6C3] = 8'h84;
mem[16'hD6C4] = 8'h20;
mem[16'hD6C5] = 8'hB1;
mem[16'hD6C6] = 8'h00;
mem[16'hD6C7] = 8'h20;
mem[16'hD6C8] = 8'h0C;
mem[16'hD6C9] = 8'hDA;
mem[16'hD6CA] = 8'hD0;
mem[16'hD6CB] = 8'hCA;
mem[16'hD6CC] = 8'h68;
mem[16'hD6CD] = 8'h68;
mem[16'hD6CE] = 8'hA5;
mem[16'hD6CF] = 8'h50;
mem[16'hD6D0] = 8'h05;
mem[16'hD6D1] = 8'h51;
mem[16'hD6D2] = 8'hD0;
mem[16'hD6D3] = 8'h06;
mem[16'hD6D4] = 8'hA9;
mem[16'hD6D5] = 8'hFF;
mem[16'hD6D6] = 8'h85;
mem[16'hD6D7] = 8'h50;
mem[16'hD6D8] = 8'h85;
mem[16'hD6D9] = 8'h51;
mem[16'hD6DA] = 8'hA0;
mem[16'hD6DB] = 8'h01;
mem[16'hD6DC] = 8'hB1;
mem[16'hD6DD] = 8'h9B;
mem[16'hD6DE] = 8'hF0;
mem[16'hD6DF] = 8'h44;
mem[16'hD6E0] = 8'h20;
mem[16'hD6E1] = 8'h58;
mem[16'hD6E2] = 8'hD8;
mem[16'hD6E3] = 8'h20;
mem[16'hD6E4] = 8'hFB;
mem[16'hD6E5] = 8'hDA;
mem[16'hD6E6] = 8'hC8;
mem[16'hD6E7] = 8'hB1;
mem[16'hD6E8] = 8'h9B;
mem[16'hD6E9] = 8'hAA;
mem[16'hD6EA] = 8'hC8;
mem[16'hD6EB] = 8'hB1;
mem[16'hD6EC] = 8'h9B;
mem[16'hD6ED] = 8'hC5;
mem[16'hD6EE] = 8'h51;
mem[16'hD6EF] = 8'hD0;
mem[16'hD6F0] = 8'h04;
mem[16'hD6F1] = 8'hE4;
mem[16'hD6F2] = 8'h50;
mem[16'hD6F3] = 8'hF0;
mem[16'hD6F4] = 8'h02;
mem[16'hD6F5] = 8'hB0;
mem[16'hD6F6] = 8'h2D;
mem[16'hD6F7] = 8'h84;
mem[16'hD6F8] = 8'h85;
mem[16'hD6F9] = 8'h20;
mem[16'hD6FA] = 8'h24;
mem[16'hD6FB] = 8'hED;
mem[16'hD6FC] = 8'hA9;
mem[16'hD6FD] = 8'h20;
mem[16'hD6FE] = 8'hA4;
mem[16'hD6FF] = 8'h85;
mem[16'hD700] = 8'h29;
mem[16'hD701] = 8'h7F;
mem[16'hD702] = 8'h20;
mem[16'hD703] = 8'h5C;
mem[16'hD704] = 8'hDB;
mem[16'hD705] = 8'hA5;
mem[16'hD706] = 8'h24;
mem[16'hD707] = 8'hC9;
mem[16'hD708] = 8'h21;
mem[16'hD709] = 8'h90;
mem[16'hD70A] = 8'h07;
mem[16'hD70B] = 8'h20;
mem[16'hD70C] = 8'hFB;
mem[16'hD70D] = 8'hDA;
mem[16'hD70E] = 8'hA9;
mem[16'hD70F] = 8'h05;
mem[16'hD710] = 8'h85;
mem[16'hD711] = 8'h24;
mem[16'hD712] = 8'hC8;
mem[16'hD713] = 8'hB1;
mem[16'hD714] = 8'h9B;
mem[16'hD715] = 8'hD0;
mem[16'hD716] = 8'h1D;
mem[16'hD717] = 8'hA8;
mem[16'hD718] = 8'hB1;
mem[16'hD719] = 8'h9B;
mem[16'hD71A] = 8'hAA;
mem[16'hD71B] = 8'hC8;
mem[16'hD71C] = 8'hB1;
mem[16'hD71D] = 8'h9B;
mem[16'hD71E] = 8'h86;
mem[16'hD71F] = 8'h9B;
mem[16'hD720] = 8'h85;
mem[16'hD721] = 8'h9C;
mem[16'hD722] = 8'hD0;
mem[16'hD723] = 8'hB6;
mem[16'hD724] = 8'hA9;
mem[16'hD725] = 8'h0D;
mem[16'hD726] = 8'h20;
mem[16'hD727] = 8'h5C;
mem[16'hD728] = 8'hDB;
mem[16'hD729] = 8'h4C;
mem[16'hD72A] = 8'hD2;
mem[16'hD72B] = 8'hD7;
mem[16'hD72C] = 8'hC8;
mem[16'hD72D] = 8'hD0;
mem[16'hD72E] = 8'h02;
mem[16'hD72F] = 8'hE6;
mem[16'hD730] = 8'h9E;
mem[16'hD731] = 8'hB1;
mem[16'hD732] = 8'h9D;
mem[16'hD733] = 8'h60;
mem[16'hD734] = 8'h10;
mem[16'hD735] = 8'hCC;
mem[16'hD736] = 8'h38;
mem[16'hD737] = 8'hE9;
mem[16'hD738] = 8'h7F;
mem[16'hD739] = 8'hAA;
mem[16'hD73A] = 8'h84;
mem[16'hD73B] = 8'h85;
mem[16'hD73C] = 8'hA0;
mem[16'hD73D] = 8'hD0;
mem[16'hD73E] = 8'h84;
mem[16'hD73F] = 8'h9D;
mem[16'hD740] = 8'hA0;
mem[16'hD741] = 8'hCF;
mem[16'hD742] = 8'h84;
mem[16'hD743] = 8'h9E;
mem[16'hD744] = 8'hA0;
mem[16'hD745] = 8'hFF;
mem[16'hD746] = 8'hCA;
mem[16'hD747] = 8'hF0;
mem[16'hD748] = 8'h07;
mem[16'hD749] = 8'h20;
mem[16'hD74A] = 8'h2C;
mem[16'hD74B] = 8'hD7;
mem[16'hD74C] = 8'h10;
mem[16'hD74D] = 8'hFB;
mem[16'hD74E] = 8'h30;
mem[16'hD74F] = 8'hF6;
mem[16'hD750] = 8'hA9;
mem[16'hD751] = 8'h20;
mem[16'hD752] = 8'h20;
mem[16'hD753] = 8'h5C;
mem[16'hD754] = 8'hDB;
mem[16'hD755] = 8'h20;
mem[16'hD756] = 8'h2C;
mem[16'hD757] = 8'hD7;
mem[16'hD758] = 8'h30;
mem[16'hD759] = 8'h05;
mem[16'hD75A] = 8'h20;
mem[16'hD75B] = 8'h5C;
mem[16'hD75C] = 8'hDB;
mem[16'hD75D] = 8'hD0;
mem[16'hD75E] = 8'hF6;
mem[16'hD75F] = 8'h20;
mem[16'hD760] = 8'h5C;
mem[16'hD761] = 8'hDB;
mem[16'hD762] = 8'hA9;
mem[16'hD763] = 8'h20;
mem[16'hD764] = 8'hD0;
mem[16'hD765] = 8'h98;
mem[16'hD766] = 8'hA9;
mem[16'hD767] = 8'h80;
mem[16'hD768] = 8'h85;
mem[16'hD769] = 8'h14;
mem[16'hD76A] = 8'h20;
mem[16'hD76B] = 8'h46;
mem[16'hD76C] = 8'hDA;
mem[16'hD76D] = 8'h20;
mem[16'hD76E] = 8'h65;
mem[16'hD76F] = 8'hD3;
mem[16'hD770] = 8'hD0;
mem[16'hD771] = 8'h05;
mem[16'hD772] = 8'h8A;
mem[16'hD773] = 8'h69;
mem[16'hD774] = 8'h0F;
mem[16'hD775] = 8'hAA;
mem[16'hD776] = 8'h9A;
mem[16'hD777] = 8'h68;
mem[16'hD778] = 8'h68;
mem[16'hD779] = 8'hA9;
mem[16'hD77A] = 8'h09;
mem[16'hD77B] = 8'h20;
mem[16'hD77C] = 8'hD6;
mem[16'hD77D] = 8'hD3;
mem[16'hD77E] = 8'h20;
mem[16'hD77F] = 8'hA3;
mem[16'hD780] = 8'hD9;
mem[16'hD781] = 8'h18;
mem[16'hD782] = 8'h98;
mem[16'hD783] = 8'h65;
mem[16'hD784] = 8'hB8;
mem[16'hD785] = 8'h48;
mem[16'hD786] = 8'hA5;
mem[16'hD787] = 8'hB9;
mem[16'hD788] = 8'h69;
mem[16'hD789] = 8'h00;
mem[16'hD78A] = 8'h48;
mem[16'hD78B] = 8'hA5;
mem[16'hD78C] = 8'h76;
mem[16'hD78D] = 8'h48;
mem[16'hD78E] = 8'hA5;
mem[16'hD78F] = 8'h75;
mem[16'hD790] = 8'h48;
mem[16'hD791] = 8'hA9;
mem[16'hD792] = 8'hC1;
mem[16'hD793] = 8'h20;
mem[16'hD794] = 8'hC0;
mem[16'hD795] = 8'hDE;
mem[16'hD796] = 8'h20;
mem[16'hD797] = 8'h6A;
mem[16'hD798] = 8'hDD;
mem[16'hD799] = 8'h20;
mem[16'hD79A] = 8'h67;
mem[16'hD79B] = 8'hDD;
mem[16'hD79C] = 8'hA5;
mem[16'hD79D] = 8'hA2;
mem[16'hD79E] = 8'h09;
mem[16'hD79F] = 8'h7F;
mem[16'hD7A0] = 8'h25;
mem[16'hD7A1] = 8'h9E;
mem[16'hD7A2] = 8'h85;
mem[16'hD7A3] = 8'h9E;
mem[16'hD7A4] = 8'hA9;
mem[16'hD7A5] = 8'hAF;
mem[16'hD7A6] = 8'hA0;
mem[16'hD7A7] = 8'hD7;
mem[16'hD7A8] = 8'h85;
mem[16'hD7A9] = 8'h5E;
mem[16'hD7AA] = 8'h84;
mem[16'hD7AB] = 8'h5F;
mem[16'hD7AC] = 8'h4C;
mem[16'hD7AD] = 8'h20;
mem[16'hD7AE] = 8'hDE;
mem[16'hD7AF] = 8'hA9;
mem[16'hD7B0] = 8'h13;
mem[16'hD7B1] = 8'hA0;
mem[16'hD7B2] = 8'hE9;
mem[16'hD7B3] = 8'h20;
mem[16'hD7B4] = 8'hF9;
mem[16'hD7B5] = 8'hEA;
mem[16'hD7B6] = 8'h20;
mem[16'hD7B7] = 8'hB7;
mem[16'hD7B8] = 8'h00;
mem[16'hD7B9] = 8'hC9;
mem[16'hD7BA] = 8'hC7;
mem[16'hD7BB] = 8'hD0;
mem[16'hD7BC] = 8'h06;
mem[16'hD7BD] = 8'h20;
mem[16'hD7BE] = 8'hB1;
mem[16'hD7BF] = 8'h00;
mem[16'hD7C0] = 8'h20;
mem[16'hD7C1] = 8'h67;
mem[16'hD7C2] = 8'hDD;
mem[16'hD7C3] = 8'h20;
mem[16'hD7C4] = 8'h82;
mem[16'hD7C5] = 8'hEB;
mem[16'hD7C6] = 8'h20;
mem[16'hD7C7] = 8'h15;
mem[16'hD7C8] = 8'hDE;
mem[16'hD7C9] = 8'hA5;
mem[16'hD7CA] = 8'h86;
mem[16'hD7CB] = 8'h48;
mem[16'hD7CC] = 8'hA5;
mem[16'hD7CD] = 8'h85;
mem[16'hD7CE] = 8'h48;
mem[16'hD7CF] = 8'hA9;
mem[16'hD7D0] = 8'h81;
mem[16'hD7D1] = 8'h48;
mem[16'hD7D2] = 8'hBA;
mem[16'hD7D3] = 8'h86;
mem[16'hD7D4] = 8'hF8;
mem[16'hD7D5] = 8'h20;
mem[16'hD7D6] = 8'h58;
mem[16'hD7D7] = 8'hD8;
mem[16'hD7D8] = 8'hA5;
mem[16'hD7D9] = 8'hB8;
mem[16'hD7DA] = 8'hA4;
mem[16'hD7DB] = 8'hB9;
mem[16'hD7DC] = 8'hA6;
mem[16'hD7DD] = 8'h76;
mem[16'hD7DE] = 8'hE8;
mem[16'hD7DF] = 8'hF0;
mem[16'hD7E0] = 8'h04;
mem[16'hD7E1] = 8'h85;
mem[16'hD7E2] = 8'h79;
mem[16'hD7E3] = 8'h84;
mem[16'hD7E4] = 8'h7A;
mem[16'hD7E5] = 8'hA0;
mem[16'hD7E6] = 8'h00;
mem[16'hD7E7] = 8'hB1;
mem[16'hD7E8] = 8'hB8;
mem[16'hD7E9] = 8'hD0;
mem[16'hD7EA] = 8'h57;
mem[16'hD7EB] = 8'hA0;
mem[16'hD7EC] = 8'h02;
mem[16'hD7ED] = 8'hB1;
mem[16'hD7EE] = 8'hB8;
mem[16'hD7EF] = 8'h18;
mem[16'hD7F0] = 8'hF0;
mem[16'hD7F1] = 8'h34;
mem[16'hD7F2] = 8'hC8;
mem[16'hD7F3] = 8'hB1;
mem[16'hD7F4] = 8'hB8;
mem[16'hD7F5] = 8'h85;
mem[16'hD7F6] = 8'h75;
mem[16'hD7F7] = 8'hC8;
mem[16'hD7F8] = 8'hB1;
mem[16'hD7F9] = 8'hB8;
mem[16'hD7FA] = 8'h85;
mem[16'hD7FB] = 8'h76;
mem[16'hD7FC] = 8'h98;
mem[16'hD7FD] = 8'h65;
mem[16'hD7FE] = 8'hB8;
mem[16'hD7FF] = 8'h85;
mem[16'hD800] = 8'hB8;
mem[16'hD801] = 8'h90;
mem[16'hD802] = 8'h02;
mem[16'hD803] = 8'hE6;
mem[16'hD804] = 8'hB9;
mem[16'hD805] = 8'h24;
mem[16'hD806] = 8'hF2;
mem[16'hD807] = 8'h10;
mem[16'hD808] = 8'h14;
mem[16'hD809] = 8'hA6;
mem[16'hD80A] = 8'h76;
mem[16'hD80B] = 8'hE8;
mem[16'hD80C] = 8'hF0;
mem[16'hD80D] = 8'h0F;
mem[16'hD80E] = 8'hA9;
mem[16'hD80F] = 8'h23;
mem[16'hD810] = 8'h20;
mem[16'hD811] = 8'h5C;
mem[16'hD812] = 8'hDB;
mem[16'hD813] = 8'hA6;
mem[16'hD814] = 8'h75;
mem[16'hD815] = 8'hA5;
mem[16'hD816] = 8'h76;
mem[16'hD817] = 8'h20;
mem[16'hD818] = 8'h24;
mem[16'hD819] = 8'hED;
mem[16'hD81A] = 8'h20;
mem[16'hD81B] = 8'h57;
mem[16'hD81C] = 8'hDB;
mem[16'hD81D] = 8'h20;
mem[16'hD81E] = 8'hB1;
mem[16'hD81F] = 8'h00;
mem[16'hD820] = 8'h20;
mem[16'hD821] = 8'h28;
mem[16'hD822] = 8'hD8;
mem[16'hD823] = 8'h4C;
mem[16'hD824] = 8'hD2;
mem[16'hD825] = 8'hD7;
mem[16'hD826] = 8'hF0;
mem[16'hD827] = 8'h62;
mem[16'hD828] = 8'hF0;
mem[16'hD829] = 8'h2D;
mem[16'hD82A] = 8'hE9;
mem[16'hD82B] = 8'h80;
mem[16'hD82C] = 8'h90;
mem[16'hD82D] = 8'h11;
mem[16'hD82E] = 8'hC9;
mem[16'hD82F] = 8'h40;
mem[16'hD830] = 8'hB0;
mem[16'hD831] = 8'h14;
mem[16'hD832] = 8'h0A;
mem[16'hD833] = 8'hA8;
mem[16'hD834] = 8'hB9;
mem[16'hD835] = 8'h01;
mem[16'hD836] = 8'hD0;
mem[16'hD837] = 8'h48;
mem[16'hD838] = 8'hB9;
mem[16'hD839] = 8'h00;
mem[16'hD83A] = 8'hD0;
mem[16'hD83B] = 8'h48;
mem[16'hD83C] = 8'h4C;
mem[16'hD83D] = 8'hB1;
mem[16'hD83E] = 8'h00;
mem[16'hD83F] = 8'h4C;
mem[16'hD840] = 8'h46;
mem[16'hD841] = 8'hDA;
mem[16'hD842] = 8'hC9;
mem[16'hD843] = 8'h3A;
mem[16'hD844] = 8'hF0;
mem[16'hD845] = 8'hBF;
mem[16'hD846] = 8'h4C;
mem[16'hD847] = 8'hC9;
mem[16'hD848] = 8'hDE;
mem[16'hD849] = 8'h38;
mem[16'hD84A] = 8'hA5;
mem[16'hD84B] = 8'h67;
mem[16'hD84C] = 8'hE9;
mem[16'hD84D] = 8'h01;
mem[16'hD84E] = 8'hA4;
mem[16'hD84F] = 8'h68;
mem[16'hD850] = 8'hB0;
mem[16'hD851] = 8'h01;
mem[16'hD852] = 8'h88;
mem[16'hD853] = 8'h85;
mem[16'hD854] = 8'h7D;
mem[16'hD855] = 8'h84;
mem[16'hD856] = 8'h7E;
mem[16'hD857] = 8'h60;
mem[16'hD858] = 8'hAD;
mem[16'hD859] = 8'h00;
mem[16'hD85A] = 8'hC0;
mem[16'hD85B] = 8'hC9;
mem[16'hD85C] = 8'h83;
mem[16'hD85D] = 8'hF0;
mem[16'hD85E] = 8'h01;
mem[16'hD85F] = 8'h60;
mem[16'hD860] = 8'h20;
mem[16'hD861] = 8'h53;
mem[16'hD862] = 8'hD5;
mem[16'hD863] = 8'hA2;
mem[16'hD864] = 8'hFF;
mem[16'hD865] = 8'h24;
mem[16'hD866] = 8'hD8;
mem[16'hD867] = 8'h10;
mem[16'hD868] = 8'h03;
mem[16'hD869] = 8'h4C;
mem[16'hD86A] = 8'hE9;
mem[16'hD86B] = 8'hF2;
mem[16'hD86C] = 8'hC9;
mem[16'hD86D] = 8'h03;
mem[16'hD86E] = 8'hB0;
mem[16'hD86F] = 8'h01;
mem[16'hD870] = 8'h18;
mem[16'hD871] = 8'hD0;
mem[16'hD872] = 8'h3C;
mem[16'hD873] = 8'hA5;
mem[16'hD874] = 8'hB8;
mem[16'hD875] = 8'hA4;
mem[16'hD876] = 8'hB9;
mem[16'hD877] = 8'hA6;
mem[16'hD878] = 8'h76;
mem[16'hD879] = 8'hE8;
mem[16'hD87A] = 8'hF0;
mem[16'hD87B] = 8'h0C;
mem[16'hD87C] = 8'h85;
mem[16'hD87D] = 8'h79;
mem[16'hD87E] = 8'h84;
mem[16'hD87F] = 8'h7A;
mem[16'hD880] = 8'hA5;
mem[16'hD881] = 8'h75;
mem[16'hD882] = 8'hA4;
mem[16'hD883] = 8'h76;
mem[16'hD884] = 8'h85;
mem[16'hD885] = 8'h77;
mem[16'hD886] = 8'h84;
mem[16'hD887] = 8'h78;
mem[16'hD888] = 8'h68;
mem[16'hD889] = 8'h68;
mem[16'hD88A] = 8'hA9;
mem[16'hD88B] = 8'h5D;
mem[16'hD88C] = 8'hA0;
mem[16'hD88D] = 8'hD3;
mem[16'hD88E] = 8'h90;
mem[16'hD88F] = 8'h03;
mem[16'hD890] = 8'h4C;
mem[16'hD891] = 8'h31;
mem[16'hD892] = 8'hD4;
mem[16'hD893] = 8'h4C;
mem[16'hD894] = 8'h3C;
mem[16'hD895] = 8'hD4;
mem[16'hD896] = 8'hD0;
mem[16'hD897] = 8'h17;
mem[16'hD898] = 8'hA2;
mem[16'hD899] = 8'hD2;
mem[16'hD89A] = 8'hA4;
mem[16'hD89B] = 8'h7A;
mem[16'hD89C] = 8'hD0;
mem[16'hD89D] = 8'h03;
mem[16'hD89E] = 8'h4C;
mem[16'hD89F] = 8'h12;
mem[16'hD8A0] = 8'hD4;
mem[16'hD8A1] = 8'hA5;
mem[16'hD8A2] = 8'h79;
mem[16'hD8A3] = 8'h85;
mem[16'hD8A4] = 8'hB8;
mem[16'hD8A5] = 8'h84;
mem[16'hD8A6] = 8'hB9;
mem[16'hD8A7] = 8'hA5;
mem[16'hD8A8] = 8'h77;
mem[16'hD8A9] = 8'hA4;
mem[16'hD8AA] = 8'h78;
mem[16'hD8AB] = 8'h85;
mem[16'hD8AC] = 8'h75;
mem[16'hD8AD] = 8'h84;
mem[16'hD8AE] = 8'h76;
mem[16'hD8AF] = 8'h60;
mem[16'hD8B0] = 8'h38;
mem[16'hD8B1] = 8'hA5;
mem[16'hD8B2] = 8'hAF;
mem[16'hD8B3] = 8'hE5;
mem[16'hD8B4] = 8'h67;
mem[16'hD8B5] = 8'h85;
mem[16'hD8B6] = 8'h50;
mem[16'hD8B7] = 8'hA5;
mem[16'hD8B8] = 8'hB0;
mem[16'hD8B9] = 8'hE5;
mem[16'hD8BA] = 8'h68;
mem[16'hD8BB] = 8'h85;
mem[16'hD8BC] = 8'h51;
mem[16'hD8BD] = 8'h20;
mem[16'hD8BE] = 8'hF0;
mem[16'hD8BF] = 8'hD8;
mem[16'hD8C0] = 8'h20;
mem[16'hD8C1] = 8'hCD;
mem[16'hD8C2] = 8'hFE;
mem[16'hD8C3] = 8'h20;
mem[16'hD8C4] = 8'h01;
mem[16'hD8C5] = 8'hD9;
mem[16'hD8C6] = 8'h4C;
mem[16'hD8C7] = 8'hCD;
mem[16'hD8C8] = 8'hFE;
mem[16'hD8C9] = 8'h20;
mem[16'hD8CA] = 8'hF0;
mem[16'hD8CB] = 8'hD8;
mem[16'hD8CC] = 8'h20;
mem[16'hD8CD] = 8'hFD;
mem[16'hD8CE] = 8'hFE;
mem[16'hD8CF] = 8'h18;
mem[16'hD8D0] = 8'hA5;
mem[16'hD8D1] = 8'h67;
mem[16'hD8D2] = 8'h65;
mem[16'hD8D3] = 8'h50;
mem[16'hD8D4] = 8'h85;
mem[16'hD8D5] = 8'h69;
mem[16'hD8D6] = 8'hA5;
mem[16'hD8D7] = 8'h68;
mem[16'hD8D8] = 8'h65;
mem[16'hD8D9] = 8'h51;
mem[16'hD8DA] = 8'h85;
mem[16'hD8DB] = 8'h6A;
mem[16'hD8DC] = 8'hA5;
mem[16'hD8DD] = 8'h52;
mem[16'hD8DE] = 8'h85;
mem[16'hD8DF] = 8'hD6;
mem[16'hD8E0] = 8'h20;
mem[16'hD8E1] = 8'h01;
mem[16'hD8E2] = 8'hD9;
mem[16'hD8E3] = 8'h20;
mem[16'hD8E4] = 8'hFD;
mem[16'hD8E5] = 8'hFE;
mem[16'hD8E6] = 8'h24;
mem[16'hD8E7] = 8'hD6;
mem[16'hD8E8] = 8'h10;
mem[16'hD8E9] = 8'h03;
mem[16'hD8EA] = 8'h4C;
mem[16'hD8EB] = 8'h65;
mem[16'hD8EC] = 8'hD6;
mem[16'hD8ED] = 8'h4C;
mem[16'hD8EE] = 8'hF2;
mem[16'hD8EF] = 8'hD4;
mem[16'hD8F0] = 8'hA9;
mem[16'hD8F1] = 8'h50;
mem[16'hD8F2] = 8'hA0;
mem[16'hD8F3] = 8'h00;
mem[16'hD8F4] = 8'h85;
mem[16'hD8F5] = 8'h3C;
mem[16'hD8F6] = 8'h84;
mem[16'hD8F7] = 8'h3D;
mem[16'hD8F8] = 8'hA9;
mem[16'hD8F9] = 8'h52;
mem[16'hD8FA] = 8'h85;
mem[16'hD8FB] = 8'h3E;
mem[16'hD8FC] = 8'h84;
mem[16'hD8FD] = 8'h3F;
mem[16'hD8FE] = 8'h84;
mem[16'hD8FF] = 8'hD6;
mem[16'hD900] = 8'h60;
mem[16'hD901] = 8'hA5;
mem[16'hD902] = 8'h67;
mem[16'hD903] = 8'hA4;
mem[16'hD904] = 8'h68;
mem[16'hD905] = 8'h85;
mem[16'hD906] = 8'h3C;
mem[16'hD907] = 8'h84;
mem[16'hD908] = 8'h3D;
mem[16'hD909] = 8'hA5;
mem[16'hD90A] = 8'h69;
mem[16'hD90B] = 8'hA4;
mem[16'hD90C] = 8'h6A;
mem[16'hD90D] = 8'h85;
mem[16'hD90E] = 8'h3E;
mem[16'hD90F] = 8'h84;
mem[16'hD910] = 8'h3F;
mem[16'hD911] = 8'h60;
mem[16'hD912] = 8'h08;
mem[16'hD913] = 8'hC6;
mem[16'hD914] = 8'h76;
mem[16'hD915] = 8'h28;
mem[16'hD916] = 8'hD0;
mem[16'hD917] = 8'h03;
mem[16'hD918] = 8'h4C;
mem[16'hD919] = 8'h65;
mem[16'hD91A] = 8'hD6;
mem[16'hD91B] = 8'h20;
mem[16'hD91C] = 8'h6C;
mem[16'hD91D] = 8'hD6;
mem[16'hD91E] = 8'h4C;
mem[16'hD91F] = 8'h35;
mem[16'hD920] = 8'hD9;
mem[16'hD921] = 8'hA9;
mem[16'hD922] = 8'h03;
mem[16'hD923] = 8'h20;
mem[16'hD924] = 8'hD6;
mem[16'hD925] = 8'hD3;
mem[16'hD926] = 8'hA5;
mem[16'hD927] = 8'hB9;
mem[16'hD928] = 8'h48;
mem[16'hD929] = 8'hA5;
mem[16'hD92A] = 8'hB8;
mem[16'hD92B] = 8'h48;
mem[16'hD92C] = 8'hA5;
mem[16'hD92D] = 8'h76;
mem[16'hD92E] = 8'h48;
mem[16'hD92F] = 8'hA5;
mem[16'hD930] = 8'h75;
mem[16'hD931] = 8'h48;
mem[16'hD932] = 8'hA9;
mem[16'hD933] = 8'hB0;
mem[16'hD934] = 8'h48;
mem[16'hD935] = 8'h20;
mem[16'hD936] = 8'hB7;
mem[16'hD937] = 8'h00;
mem[16'hD938] = 8'h20;
mem[16'hD939] = 8'h3E;
mem[16'hD93A] = 8'hD9;
mem[16'hD93B] = 8'h4C;
mem[16'hD93C] = 8'hD2;
mem[16'hD93D] = 8'hD7;
mem[16'hD93E] = 8'h20;
mem[16'hD93F] = 8'h0C;
mem[16'hD940] = 8'hDA;
mem[16'hD941] = 8'h20;
mem[16'hD942] = 8'hA6;
mem[16'hD943] = 8'hD9;
mem[16'hD944] = 8'hA5;
mem[16'hD945] = 8'h76;
mem[16'hD946] = 8'hC5;
mem[16'hD947] = 8'h51;
mem[16'hD948] = 8'hB0;
mem[16'hD949] = 8'h0B;
mem[16'hD94A] = 8'h98;
mem[16'hD94B] = 8'h38;
mem[16'hD94C] = 8'h65;
mem[16'hD94D] = 8'hB8;
mem[16'hD94E] = 8'hA6;
mem[16'hD94F] = 8'hB9;
mem[16'hD950] = 8'h90;
mem[16'hD951] = 8'h07;
mem[16'hD952] = 8'hE8;
mem[16'hD953] = 8'hB0;
mem[16'hD954] = 8'h04;
mem[16'hD955] = 8'hA5;
mem[16'hD956] = 8'h67;
mem[16'hD957] = 8'hA6;
mem[16'hD958] = 8'h68;
mem[16'hD959] = 8'h20;
mem[16'hD95A] = 8'h1E;
mem[16'hD95B] = 8'hD6;
mem[16'hD95C] = 8'h90;
mem[16'hD95D] = 8'h1E;
mem[16'hD95E] = 8'hA5;
mem[16'hD95F] = 8'h9B;
mem[16'hD960] = 8'hE9;
mem[16'hD961] = 8'h01;
mem[16'hD962] = 8'h85;
mem[16'hD963] = 8'hB8;
mem[16'hD964] = 8'hA5;
mem[16'hD965] = 8'h9C;
mem[16'hD966] = 8'hE9;
mem[16'hD967] = 8'h00;
mem[16'hD968] = 8'h85;
mem[16'hD969] = 8'hB9;
mem[16'hD96A] = 8'h60;
mem[16'hD96B] = 8'hD0;
mem[16'hD96C] = 8'hFD;
mem[16'hD96D] = 8'hA9;
mem[16'hD96E] = 8'hFF;
mem[16'hD96F] = 8'h85;
mem[16'hD970] = 8'h85;
mem[16'hD971] = 8'h20;
mem[16'hD972] = 8'h65;
mem[16'hD973] = 8'hD3;
mem[16'hD974] = 8'h9A;
mem[16'hD975] = 8'hC9;
mem[16'hD976] = 8'hB0;
mem[16'hD977] = 8'hF0;
mem[16'hD978] = 8'h0B;
mem[16'hD979] = 8'hA2;
mem[16'hD97A] = 8'h16;
mem[16'hD97B] = 8'h2C;
mem[16'hD97C] = 8'hA2;
mem[16'hD97D] = 8'h5A;
mem[16'hD97E] = 8'h4C;
mem[16'hD97F] = 8'h12;
mem[16'hD980] = 8'hD4;
mem[16'hD981] = 8'h4C;
mem[16'hD982] = 8'hC9;
mem[16'hD983] = 8'hDE;
mem[16'hD984] = 8'h68;
mem[16'hD985] = 8'h68;
mem[16'hD986] = 8'hC0;
mem[16'hD987] = 8'h42;
mem[16'hD988] = 8'hF0;
mem[16'hD989] = 8'h3B;
mem[16'hD98A] = 8'h85;
mem[16'hD98B] = 8'h75;
mem[16'hD98C] = 8'h68;
mem[16'hD98D] = 8'h85;
mem[16'hD98E] = 8'h76;
mem[16'hD98F] = 8'h68;
mem[16'hD990] = 8'h85;
mem[16'hD991] = 8'hB8;
mem[16'hD992] = 8'h68;
mem[16'hD993] = 8'h85;
mem[16'hD994] = 8'hB9;
mem[16'hD995] = 8'h20;
mem[16'hD996] = 8'hA3;
mem[16'hD997] = 8'hD9;
mem[16'hD998] = 8'h98;
mem[16'hD999] = 8'h18;
mem[16'hD99A] = 8'h65;
mem[16'hD99B] = 8'hB8;
mem[16'hD99C] = 8'h85;
mem[16'hD99D] = 8'hB8;
mem[16'hD99E] = 8'h90;
mem[16'hD99F] = 8'h02;
mem[16'hD9A0] = 8'hE6;
mem[16'hD9A1] = 8'hB9;
mem[16'hD9A2] = 8'h60;
mem[16'hD9A3] = 8'hA2;
mem[16'hD9A4] = 8'h3A;
mem[16'hD9A5] = 8'h2C;
mem[16'hD9A6] = 8'hA2;
mem[16'hD9A7] = 8'h00;
mem[16'hD9A8] = 8'h86;
mem[16'hD9A9] = 8'h0D;
mem[16'hD9AA] = 8'hA0;
mem[16'hD9AB] = 8'h00;
mem[16'hD9AC] = 8'h84;
mem[16'hD9AD] = 8'h0E;
mem[16'hD9AE] = 8'hA5;
mem[16'hD9AF] = 8'h0E;
mem[16'hD9B0] = 8'hA6;
mem[16'hD9B1] = 8'h0D;
mem[16'hD9B2] = 8'h85;
mem[16'hD9B3] = 8'h0D;
mem[16'hD9B4] = 8'h86;
mem[16'hD9B5] = 8'h0E;
mem[16'hD9B6] = 8'hB1;
mem[16'hD9B7] = 8'hB8;
mem[16'hD9B8] = 8'hF0;
mem[16'hD9B9] = 8'hE8;
mem[16'hD9BA] = 8'hC5;
mem[16'hD9BB] = 8'h0E;
mem[16'hD9BC] = 8'hF0;
mem[16'hD9BD] = 8'hE4;
mem[16'hD9BE] = 8'hC8;
mem[16'hD9BF] = 8'hC9;
mem[16'hD9C0] = 8'h22;
mem[16'hD9C1] = 8'hD0;
mem[16'hD9C2] = 8'hF3;
mem[16'hD9C3] = 8'hF0;
mem[16'hD9C4] = 8'hE9;
mem[16'hD9C5] = 8'h68;
mem[16'hD9C6] = 8'h68;
mem[16'hD9C7] = 8'h68;
mem[16'hD9C8] = 8'h60;
mem[16'hD9C9] = 8'h20;
mem[16'hD9CA] = 8'h7B;
mem[16'hD9CB] = 8'hDD;
mem[16'hD9CC] = 8'h20;
mem[16'hD9CD] = 8'hB7;
mem[16'hD9CE] = 8'h00;
mem[16'hD9CF] = 8'hC9;
mem[16'hD9D0] = 8'hAB;
mem[16'hD9D1] = 8'hF0;
mem[16'hD9D2] = 8'h05;
mem[16'hD9D3] = 8'hA9;
mem[16'hD9D4] = 8'hC4;
mem[16'hD9D5] = 8'h20;
mem[16'hD9D6] = 8'hC0;
mem[16'hD9D7] = 8'hDE;
mem[16'hD9D8] = 8'hA5;
mem[16'hD9D9] = 8'h9D;
mem[16'hD9DA] = 8'hD0;
mem[16'hD9DB] = 8'h05;
mem[16'hD9DC] = 8'h20;
mem[16'hD9DD] = 8'hA6;
mem[16'hD9DE] = 8'hD9;
mem[16'hD9DF] = 8'hF0;
mem[16'hD9E0] = 8'hB7;
mem[16'hD9E1] = 8'h20;
mem[16'hD9E2] = 8'hB7;
mem[16'hD9E3] = 8'h00;
mem[16'hD9E4] = 8'hB0;
mem[16'hD9E5] = 8'h03;
mem[16'hD9E6] = 8'h4C;
mem[16'hD9E7] = 8'h3E;
mem[16'hD9E8] = 8'hD9;
mem[16'hD9E9] = 8'h4C;
mem[16'hD9EA] = 8'h28;
mem[16'hD9EB] = 8'hD8;
mem[16'hD9EC] = 8'h20;
mem[16'hD9ED] = 8'hF8;
mem[16'hD9EE] = 8'hE6;
mem[16'hD9EF] = 8'h48;
mem[16'hD9F0] = 8'hC9;
mem[16'hD9F1] = 8'hB0;
mem[16'hD9F2] = 8'hF0;
mem[16'hD9F3] = 8'h04;
mem[16'hD9F4] = 8'hC9;
mem[16'hD9F5] = 8'hAB;
mem[16'hD9F6] = 8'hD0;
mem[16'hD9F7] = 8'h89;
mem[16'hD9F8] = 8'hC6;
mem[16'hD9F9] = 8'hA1;
mem[16'hD9FA] = 8'hD0;
mem[16'hD9FB] = 8'h04;
mem[16'hD9FC] = 8'h68;
mem[16'hD9FD] = 8'h4C;
mem[16'hD9FE] = 8'h2A;
mem[16'hD9FF] = 8'hD8;
mem[16'hDA00] = 8'h20;
mem[16'hDA01] = 8'hB1;
mem[16'hDA02] = 8'h00;
mem[16'hDA03] = 8'h20;
mem[16'hDA04] = 8'h0C;
mem[16'hDA05] = 8'hDA;
mem[16'hDA06] = 8'hC9;
mem[16'hDA07] = 8'h2C;
mem[16'hDA08] = 8'hF0;
mem[16'hDA09] = 8'hEE;
mem[16'hDA0A] = 8'h68;
mem[16'hDA0B] = 8'h60;
mem[16'hDA0C] = 8'hA2;
mem[16'hDA0D] = 8'h00;
mem[16'hDA0E] = 8'h86;
mem[16'hDA0F] = 8'h50;
mem[16'hDA10] = 8'h86;
mem[16'hDA11] = 8'h51;
mem[16'hDA12] = 8'hB0;
mem[16'hDA13] = 8'hF7;
mem[16'hDA14] = 8'hE9;
mem[16'hDA15] = 8'h2F;
mem[16'hDA16] = 8'h85;
mem[16'hDA17] = 8'h0D;
mem[16'hDA18] = 8'hA5;
mem[16'hDA19] = 8'h51;
mem[16'hDA1A] = 8'h85;
mem[16'hDA1B] = 8'h5E;
mem[16'hDA1C] = 8'hC9;
mem[16'hDA1D] = 8'h19;
mem[16'hDA1E] = 8'hB0;
mem[16'hDA1F] = 8'hD4;
mem[16'hDA20] = 8'hA5;
mem[16'hDA21] = 8'h50;
mem[16'hDA22] = 8'h0A;
mem[16'hDA23] = 8'h26;
mem[16'hDA24] = 8'h5E;
mem[16'hDA25] = 8'h0A;
mem[16'hDA26] = 8'h26;
mem[16'hDA27] = 8'h5E;
mem[16'hDA28] = 8'h65;
mem[16'hDA29] = 8'h50;
mem[16'hDA2A] = 8'h85;
mem[16'hDA2B] = 8'h50;
mem[16'hDA2C] = 8'hA5;
mem[16'hDA2D] = 8'h5E;
mem[16'hDA2E] = 8'h65;
mem[16'hDA2F] = 8'h51;
mem[16'hDA30] = 8'h85;
mem[16'hDA31] = 8'h51;
mem[16'hDA32] = 8'h06;
mem[16'hDA33] = 8'h50;
mem[16'hDA34] = 8'h26;
mem[16'hDA35] = 8'h51;
mem[16'hDA36] = 8'hA5;
mem[16'hDA37] = 8'h50;
mem[16'hDA38] = 8'h65;
mem[16'hDA39] = 8'h0D;
mem[16'hDA3A] = 8'h85;
mem[16'hDA3B] = 8'h50;
mem[16'hDA3C] = 8'h90;
mem[16'hDA3D] = 8'h02;
mem[16'hDA3E] = 8'hE6;
mem[16'hDA3F] = 8'h51;
mem[16'hDA40] = 8'h20;
mem[16'hDA41] = 8'hB1;
mem[16'hDA42] = 8'h00;
mem[16'hDA43] = 8'h4C;
mem[16'hDA44] = 8'h12;
mem[16'hDA45] = 8'hDA;
mem[16'hDA46] = 8'h20;
mem[16'hDA47] = 8'hE3;
mem[16'hDA48] = 8'hDF;
mem[16'hDA49] = 8'h85;
mem[16'hDA4A] = 8'h85;
mem[16'hDA4B] = 8'h84;
mem[16'hDA4C] = 8'h86;
mem[16'hDA4D] = 8'hA9;
mem[16'hDA4E] = 8'hD0;
mem[16'hDA4F] = 8'h20;
mem[16'hDA50] = 8'hC0;
mem[16'hDA51] = 8'hDE;
mem[16'hDA52] = 8'hA5;
mem[16'hDA53] = 8'h12;
mem[16'hDA54] = 8'h48;
mem[16'hDA55] = 8'hA5;
mem[16'hDA56] = 8'h11;
mem[16'hDA57] = 8'h48;
mem[16'hDA58] = 8'h20;
mem[16'hDA59] = 8'h7B;
mem[16'hDA5A] = 8'hDD;
mem[16'hDA5B] = 8'h68;
mem[16'hDA5C] = 8'h2A;
mem[16'hDA5D] = 8'h20;
mem[16'hDA5E] = 8'h6D;
mem[16'hDA5F] = 8'hDD;
mem[16'hDA60] = 8'hD0;
mem[16'hDA61] = 8'h18;
mem[16'hDA62] = 8'h68;
mem[16'hDA63] = 8'h10;
mem[16'hDA64] = 8'h12;
mem[16'hDA65] = 8'h20;
mem[16'hDA66] = 8'h72;
mem[16'hDA67] = 8'hEB;
mem[16'hDA68] = 8'h20;
mem[16'hDA69] = 8'h0C;
mem[16'hDA6A] = 8'hE1;
mem[16'hDA6B] = 8'hA0;
mem[16'hDA6C] = 8'h00;
mem[16'hDA6D] = 8'hA5;
mem[16'hDA6E] = 8'hA0;
mem[16'hDA6F] = 8'h91;
mem[16'hDA70] = 8'h85;
mem[16'hDA71] = 8'hC8;
mem[16'hDA72] = 8'hA5;
mem[16'hDA73] = 8'hA1;
mem[16'hDA74] = 8'h91;
mem[16'hDA75] = 8'h85;
mem[16'hDA76] = 8'h60;
mem[16'hDA77] = 8'h4C;
mem[16'hDA78] = 8'h27;
mem[16'hDA79] = 8'hEB;
mem[16'hDA7A] = 8'h68;
mem[16'hDA7B] = 8'hA0;
mem[16'hDA7C] = 8'h02;
mem[16'hDA7D] = 8'hB1;
mem[16'hDA7E] = 8'hA0;
mem[16'hDA7F] = 8'hC5;
mem[16'hDA80] = 8'h70;
mem[16'hDA81] = 8'h90;
mem[16'hDA82] = 8'h17;
mem[16'hDA83] = 8'hD0;
mem[16'hDA84] = 8'h07;
mem[16'hDA85] = 8'h88;
mem[16'hDA86] = 8'hB1;
mem[16'hDA87] = 8'hA0;
mem[16'hDA88] = 8'hC5;
mem[16'hDA89] = 8'h6F;
mem[16'hDA8A] = 8'h90;
mem[16'hDA8B] = 8'h0E;
mem[16'hDA8C] = 8'hA4;
mem[16'hDA8D] = 8'hA1;
mem[16'hDA8E] = 8'hC4;
mem[16'hDA8F] = 8'h6A;
mem[16'hDA90] = 8'h90;
mem[16'hDA91] = 8'h08;
mem[16'hDA92] = 8'hD0;
mem[16'hDA93] = 8'h0D;
mem[16'hDA94] = 8'hA5;
mem[16'hDA95] = 8'hA0;
mem[16'hDA96] = 8'hC5;
mem[16'hDA97] = 8'h69;
mem[16'hDA98] = 8'hB0;
mem[16'hDA99] = 8'h07;
mem[16'hDA9A] = 8'hA5;
mem[16'hDA9B] = 8'hA0;
mem[16'hDA9C] = 8'hA4;
mem[16'hDA9D] = 8'hA1;
mem[16'hDA9E] = 8'h4C;
mem[16'hDA9F] = 8'hB7;
mem[16'hDAA0] = 8'hDA;
mem[16'hDAA1] = 8'hA0;
mem[16'hDAA2] = 8'h00;
mem[16'hDAA3] = 8'hB1;
mem[16'hDAA4] = 8'hA0;
mem[16'hDAA5] = 8'h20;
mem[16'hDAA6] = 8'hD5;
mem[16'hDAA7] = 8'hE3;
mem[16'hDAA8] = 8'hA5;
mem[16'hDAA9] = 8'h8C;
mem[16'hDAAA] = 8'hA4;
mem[16'hDAAB] = 8'h8D;
mem[16'hDAAC] = 8'h85;
mem[16'hDAAD] = 8'hAB;
mem[16'hDAAE] = 8'h84;
mem[16'hDAAF] = 8'hAC;
mem[16'hDAB0] = 8'h20;
mem[16'hDAB1] = 8'hD4;
mem[16'hDAB2] = 8'hE5;
mem[16'hDAB3] = 8'hA9;
mem[16'hDAB4] = 8'h9D;
mem[16'hDAB5] = 8'hA0;
mem[16'hDAB6] = 8'h00;
mem[16'hDAB7] = 8'h85;
mem[16'hDAB8] = 8'h8C;
mem[16'hDAB9] = 8'h84;
mem[16'hDABA] = 8'h8D;
mem[16'hDABB] = 8'h20;
mem[16'hDABC] = 8'h35;
mem[16'hDABD] = 8'hE6;
mem[16'hDABE] = 8'hA0;
mem[16'hDABF] = 8'h00;
mem[16'hDAC0] = 8'hB1;
mem[16'hDAC1] = 8'h8C;
mem[16'hDAC2] = 8'h91;
mem[16'hDAC3] = 8'h85;
mem[16'hDAC4] = 8'hC8;
mem[16'hDAC5] = 8'hB1;
mem[16'hDAC6] = 8'h8C;
mem[16'hDAC7] = 8'h91;
mem[16'hDAC8] = 8'h85;
mem[16'hDAC9] = 8'hC8;
mem[16'hDACA] = 8'hB1;
mem[16'hDACB] = 8'h8C;
mem[16'hDACC] = 8'h91;
mem[16'hDACD] = 8'h85;
mem[16'hDACE] = 8'h60;
mem[16'hDACF] = 8'h20;
mem[16'hDAD0] = 8'h3D;
mem[16'hDAD1] = 8'hDB;
mem[16'hDAD2] = 8'h20;
mem[16'hDAD3] = 8'hB7;
mem[16'hDAD4] = 8'h00;
mem[16'hDAD5] = 8'hF0;
mem[16'hDAD6] = 8'h24;
mem[16'hDAD7] = 8'hF0;
mem[16'hDAD8] = 8'h29;
mem[16'hDAD9] = 8'hC9;
mem[16'hDADA] = 8'hC0;
mem[16'hDADB] = 8'hF0;
mem[16'hDADC] = 8'h39;
mem[16'hDADD] = 8'hC9;
mem[16'hDADE] = 8'hC3;
mem[16'hDADF] = 8'h18;
mem[16'hDAE0] = 8'hF0;
mem[16'hDAE1] = 8'h34;
mem[16'hDAE2] = 8'hC9;
mem[16'hDAE3] = 8'h2C;
mem[16'hDAE4] = 8'h18;
mem[16'hDAE5] = 8'hF0;
mem[16'hDAE6] = 8'h1C;
mem[16'hDAE7] = 8'hC9;
mem[16'hDAE8] = 8'h3B;
mem[16'hDAE9] = 8'hF0;
mem[16'hDAEA] = 8'h44;
mem[16'hDAEB] = 8'h20;
mem[16'hDAEC] = 8'h7B;
mem[16'hDAED] = 8'hDD;
mem[16'hDAEE] = 8'h24;
mem[16'hDAEF] = 8'h11;
mem[16'hDAF0] = 8'h30;
mem[16'hDAF1] = 8'hDD;
mem[16'hDAF2] = 8'h20;
mem[16'hDAF3] = 8'h34;
mem[16'hDAF4] = 8'hED;
mem[16'hDAF5] = 8'h20;
mem[16'hDAF6] = 8'hE7;
mem[16'hDAF7] = 8'hE3;
mem[16'hDAF8] = 8'h4C;
mem[16'hDAF9] = 8'hCF;
mem[16'hDAFA] = 8'hDA;
mem[16'hDAFB] = 8'hA9;
mem[16'hDAFC] = 8'h0D;
mem[16'hDAFD] = 8'h20;
mem[16'hDAFE] = 8'h5C;
mem[16'hDAFF] = 8'hDB;
mem[16'hDB00] = 8'h49;
mem[16'hDB01] = 8'hFF;
mem[16'hDB02] = 8'h60;
mem[16'hDB03] = 8'hA5;
mem[16'hDB04] = 8'h24;
mem[16'hDB05] = 8'hC9;
mem[16'hDB06] = 8'h18;
mem[16'hDB07] = 8'h90;
mem[16'hDB08] = 8'h05;
mem[16'hDB09] = 8'h20;
mem[16'hDB0A] = 8'hFB;
mem[16'hDB0B] = 8'hDA;
mem[16'hDB0C] = 8'hD0;
mem[16'hDB0D] = 8'h21;
mem[16'hDB0E] = 8'h69;
mem[16'hDB0F] = 8'h10;
mem[16'hDB10] = 8'h29;
mem[16'hDB11] = 8'hF0;
mem[16'hDB12] = 8'h85;
mem[16'hDB13] = 8'h24;
mem[16'hDB14] = 8'h90;
mem[16'hDB15] = 8'h19;
mem[16'hDB16] = 8'h08;
mem[16'hDB17] = 8'h20;
mem[16'hDB18] = 8'hF5;
mem[16'hDB19] = 8'hE6;
mem[16'hDB1A] = 8'hC9;
mem[16'hDB1B] = 8'h29;
mem[16'hDB1C] = 8'hF0;
mem[16'hDB1D] = 8'h03;
mem[16'hDB1E] = 8'h4C;
mem[16'hDB1F] = 8'hC9;
mem[16'hDB20] = 8'hDE;
mem[16'hDB21] = 8'h28;
mem[16'hDB22] = 8'h90;
mem[16'hDB23] = 8'h07;
mem[16'hDB24] = 8'hCA;
mem[16'hDB25] = 8'h8A;
mem[16'hDB26] = 8'hE5;
mem[16'hDB27] = 8'h24;
mem[16'hDB28] = 8'h90;
mem[16'hDB29] = 8'h05;
mem[16'hDB2A] = 8'hAA;
mem[16'hDB2B] = 8'hE8;
mem[16'hDB2C] = 8'hCA;
mem[16'hDB2D] = 8'hD0;
mem[16'hDB2E] = 8'h06;
mem[16'hDB2F] = 8'h20;
mem[16'hDB30] = 8'hB1;
mem[16'hDB31] = 8'h00;
mem[16'hDB32] = 8'h4C;
mem[16'hDB33] = 8'hD7;
mem[16'hDB34] = 8'hDA;
mem[16'hDB35] = 8'h20;
mem[16'hDB36] = 8'h57;
mem[16'hDB37] = 8'hDB;
mem[16'hDB38] = 8'hD0;
mem[16'hDB39] = 8'hF2;
mem[16'hDB3A] = 8'h20;
mem[16'hDB3B] = 8'hE7;
mem[16'hDB3C] = 8'hE3;
mem[16'hDB3D] = 8'h20;
mem[16'hDB3E] = 8'h00;
mem[16'hDB3F] = 8'hE6;
mem[16'hDB40] = 8'hAA;
mem[16'hDB41] = 8'hA0;
mem[16'hDB42] = 8'h00;
mem[16'hDB43] = 8'hE8;
mem[16'hDB44] = 8'hCA;
mem[16'hDB45] = 8'hF0;
mem[16'hDB46] = 8'hBB;
mem[16'hDB47] = 8'hB1;
mem[16'hDB48] = 8'h5E;
mem[16'hDB49] = 8'h20;
mem[16'hDB4A] = 8'h5C;
mem[16'hDB4B] = 8'hDB;
mem[16'hDB4C] = 8'hC8;
mem[16'hDB4D] = 8'hC9;
mem[16'hDB4E] = 8'h0D;
mem[16'hDB4F] = 8'hD0;
mem[16'hDB50] = 8'hF3;
mem[16'hDB51] = 8'h20;
mem[16'hDB52] = 8'h00;
mem[16'hDB53] = 8'hDB;
mem[16'hDB54] = 8'h4C;
mem[16'hDB55] = 8'h44;
mem[16'hDB56] = 8'hDB;
mem[16'hDB57] = 8'hA9;
mem[16'hDB58] = 8'h20;
mem[16'hDB59] = 8'h2C;
mem[16'hDB5A] = 8'hA9;
mem[16'hDB5B] = 8'h3F;
mem[16'hDB5C] = 8'h09;
mem[16'hDB5D] = 8'h80;
mem[16'hDB5E] = 8'hC9;
mem[16'hDB5F] = 8'hA0;
mem[16'hDB60] = 8'h90;
mem[16'hDB61] = 8'h02;
mem[16'hDB62] = 8'h05;
mem[16'hDB63] = 8'hF3;
mem[16'hDB64] = 8'h20;
mem[16'hDB65] = 8'hED;
mem[16'hDB66] = 8'hFD;
mem[16'hDB67] = 8'h29;
mem[16'hDB68] = 8'h7F;
mem[16'hDB69] = 8'h48;
mem[16'hDB6A] = 8'hA5;
mem[16'hDB6B] = 8'hF1;
mem[16'hDB6C] = 8'h20;
mem[16'hDB6D] = 8'hA8;
mem[16'hDB6E] = 8'hFC;
mem[16'hDB6F] = 8'h68;
mem[16'hDB70] = 8'h60;
mem[16'hDB71] = 8'hA5;
mem[16'hDB72] = 8'h15;
mem[16'hDB73] = 8'hF0;
mem[16'hDB74] = 8'h12;
mem[16'hDB75] = 8'h30;
mem[16'hDB76] = 8'h04;
mem[16'hDB77] = 8'hA0;
mem[16'hDB78] = 8'hFF;
mem[16'hDB79] = 8'hD0;
mem[16'hDB7A] = 8'h04;
mem[16'hDB7B] = 8'hA5;
mem[16'hDB7C] = 8'h7B;
mem[16'hDB7D] = 8'hA4;
mem[16'hDB7E] = 8'h7C;
mem[16'hDB7F] = 8'h85;
mem[16'hDB80] = 8'h75;
mem[16'hDB81] = 8'h84;
mem[16'hDB82] = 8'h76;
mem[16'hDB83] = 8'h4C;
mem[16'hDB84] = 8'hC9;
mem[16'hDB85] = 8'hDE;
mem[16'hDB86] = 8'h68;
mem[16'hDB87] = 8'h24;
mem[16'hDB88] = 8'hD8;
mem[16'hDB89] = 8'h10;
mem[16'hDB8A] = 8'h05;
mem[16'hDB8B] = 8'hA2;
mem[16'hDB8C] = 8'hFE;
mem[16'hDB8D] = 8'h4C;
mem[16'hDB8E] = 8'hE9;
mem[16'hDB8F] = 8'hF2;
mem[16'hDB90] = 8'hA9;
mem[16'hDB91] = 8'hEF;
mem[16'hDB92] = 8'hA0;
mem[16'hDB93] = 8'hDC;
mem[16'hDB94] = 8'h20;
mem[16'hDB95] = 8'h3A;
mem[16'hDB96] = 8'hDB;
mem[16'hDB97] = 8'hA5;
mem[16'hDB98] = 8'h79;
mem[16'hDB99] = 8'hA4;
mem[16'hDB9A] = 8'h7A;
mem[16'hDB9B] = 8'h85;
mem[16'hDB9C] = 8'hB8;
mem[16'hDB9D] = 8'h84;
mem[16'hDB9E] = 8'hB9;
mem[16'hDB9F] = 8'h60;
mem[16'hDBA0] = 8'h20;
mem[16'hDBA1] = 8'h06;
mem[16'hDBA2] = 8'hE3;
mem[16'hDBA3] = 8'hA2;
mem[16'hDBA4] = 8'h01;
mem[16'hDBA5] = 8'hA0;
mem[16'hDBA6] = 8'h02;
mem[16'hDBA7] = 8'hA9;
mem[16'hDBA8] = 8'h00;
mem[16'hDBA9] = 8'h8D;
mem[16'hDBAA] = 8'h01;
mem[16'hDBAB] = 8'h02;
mem[16'hDBAC] = 8'hA9;
mem[16'hDBAD] = 8'h40;
mem[16'hDBAE] = 8'h20;
mem[16'hDBAF] = 8'hEB;
mem[16'hDBB0] = 8'hDB;
mem[16'hDBB1] = 8'h60;
mem[16'hDBB2] = 8'hC9;
mem[16'hDBB3] = 8'h22;
mem[16'hDBB4] = 8'hD0;
mem[16'hDBB5] = 8'h0E;
mem[16'hDBB6] = 8'h20;
mem[16'hDBB7] = 8'h81;
mem[16'hDBB8] = 8'hDE;
mem[16'hDBB9] = 8'hA9;
mem[16'hDBBA] = 8'h3B;
mem[16'hDBBB] = 8'h20;
mem[16'hDBBC] = 8'hC0;
mem[16'hDBBD] = 8'hDE;
mem[16'hDBBE] = 8'h20;
mem[16'hDBBF] = 8'h3D;
mem[16'hDBC0] = 8'hDB;
mem[16'hDBC1] = 8'h4C;
mem[16'hDBC2] = 8'hC7;
mem[16'hDBC3] = 8'hDB;
mem[16'hDBC4] = 8'h20;
mem[16'hDBC5] = 8'h5A;
mem[16'hDBC6] = 8'hDB;
mem[16'hDBC7] = 8'h20;
mem[16'hDBC8] = 8'h06;
mem[16'hDBC9] = 8'hE3;
mem[16'hDBCA] = 8'hA9;
mem[16'hDBCB] = 8'h2C;
mem[16'hDBCC] = 8'h8D;
mem[16'hDBCD] = 8'hFF;
mem[16'hDBCE] = 8'h01;
mem[16'hDBCF] = 8'h20;
mem[16'hDBD0] = 8'h2C;
mem[16'hDBD1] = 8'hD5;
mem[16'hDBD2] = 8'hAD;
mem[16'hDBD3] = 8'h00;
mem[16'hDBD4] = 8'h02;
mem[16'hDBD5] = 8'hC9;
mem[16'hDBD6] = 8'h03;
mem[16'hDBD7] = 8'hD0;
mem[16'hDBD8] = 8'h10;
mem[16'hDBD9] = 8'h4C;
mem[16'hDBDA] = 8'h63;
mem[16'hDBDB] = 8'hD8;
mem[16'hDBDC] = 8'h20;
mem[16'hDBDD] = 8'h5A;
mem[16'hDBDE] = 8'hDB;
mem[16'hDBDF] = 8'h4C;
mem[16'hDBE0] = 8'h2C;
mem[16'hDBE1] = 8'hD5;
mem[16'hDBE2] = 8'hA6;
mem[16'hDBE3] = 8'h7D;
mem[16'hDBE4] = 8'hA4;
mem[16'hDBE5] = 8'h7E;
mem[16'hDBE6] = 8'hA9;
mem[16'hDBE7] = 8'h98;
mem[16'hDBE8] = 8'h2C;
mem[16'hDBE9] = 8'hA9;
mem[16'hDBEA] = 8'h00;
mem[16'hDBEB] = 8'h85;
mem[16'hDBEC] = 8'h15;
mem[16'hDBED] = 8'h86;
mem[16'hDBEE] = 8'h7F;
mem[16'hDBEF] = 8'h84;
mem[16'hDBF0] = 8'h80;
mem[16'hDBF1] = 8'h20;
mem[16'hDBF2] = 8'hE3;
mem[16'hDBF3] = 8'hDF;
mem[16'hDBF4] = 8'h85;
mem[16'hDBF5] = 8'h85;
mem[16'hDBF6] = 8'h84;
mem[16'hDBF7] = 8'h86;
mem[16'hDBF8] = 8'hA5;
mem[16'hDBF9] = 8'hB8;
mem[16'hDBFA] = 8'hA4;
mem[16'hDBFB] = 8'hB9;
mem[16'hDBFC] = 8'h85;
mem[16'hDBFD] = 8'h87;
mem[16'hDBFE] = 8'h84;
mem[16'hDBFF] = 8'h88;
mem[16'hDC00] = 8'hA6;
mem[16'hDC01] = 8'h7F;
mem[16'hDC02] = 8'hA4;
mem[16'hDC03] = 8'h80;
mem[16'hDC04] = 8'h86;
mem[16'hDC05] = 8'hB8;
mem[16'hDC06] = 8'h84;
mem[16'hDC07] = 8'hB9;
mem[16'hDC08] = 8'h20;
mem[16'hDC09] = 8'hB7;
mem[16'hDC0A] = 8'h00;
mem[16'hDC0B] = 8'hD0;
mem[16'hDC0C] = 8'h1E;
mem[16'hDC0D] = 8'h24;
mem[16'hDC0E] = 8'h15;
mem[16'hDC0F] = 8'h50;
mem[16'hDC10] = 8'h0E;
mem[16'hDC11] = 8'h20;
mem[16'hDC12] = 8'h0C;
mem[16'hDC13] = 8'hFD;
mem[16'hDC14] = 8'h29;
mem[16'hDC15] = 8'h7F;
mem[16'hDC16] = 8'h8D;
mem[16'hDC17] = 8'h00;
mem[16'hDC18] = 8'h02;
mem[16'hDC19] = 8'hA2;
mem[16'hDC1A] = 8'hFF;
mem[16'hDC1B] = 8'hA0;
mem[16'hDC1C] = 8'h01;
mem[16'hDC1D] = 8'hD0;
mem[16'hDC1E] = 8'h08;
mem[16'hDC1F] = 8'h30;
mem[16'hDC20] = 8'h7F;
mem[16'hDC21] = 8'h20;
mem[16'hDC22] = 8'h5A;
mem[16'hDC23] = 8'hDB;
mem[16'hDC24] = 8'h20;
mem[16'hDC25] = 8'hDC;
mem[16'hDC26] = 8'hDB;
mem[16'hDC27] = 8'h86;
mem[16'hDC28] = 8'hB8;
mem[16'hDC29] = 8'h84;
mem[16'hDC2A] = 8'hB9;
mem[16'hDC2B] = 8'h20;
mem[16'hDC2C] = 8'hB1;
mem[16'hDC2D] = 8'h00;
mem[16'hDC2E] = 8'h24;
mem[16'hDC2F] = 8'h11;
mem[16'hDC30] = 8'h10;
mem[16'hDC31] = 8'h31;
mem[16'hDC32] = 8'h24;
mem[16'hDC33] = 8'h15;
mem[16'hDC34] = 8'h50;
mem[16'hDC35] = 8'h09;
mem[16'hDC36] = 8'hE8;
mem[16'hDC37] = 8'h86;
mem[16'hDC38] = 8'hB8;
mem[16'hDC39] = 8'hA9;
mem[16'hDC3A] = 8'h00;
mem[16'hDC3B] = 8'h85;
mem[16'hDC3C] = 8'h0D;
mem[16'hDC3D] = 8'hF0;
mem[16'hDC3E] = 8'h0C;
mem[16'hDC3F] = 8'h85;
mem[16'hDC40] = 8'h0D;
mem[16'hDC41] = 8'hC9;
mem[16'hDC42] = 8'h22;
mem[16'hDC43] = 8'hF0;
mem[16'hDC44] = 8'h07;
mem[16'hDC45] = 8'hA9;
mem[16'hDC46] = 8'h3A;
mem[16'hDC47] = 8'h85;
mem[16'hDC48] = 8'h0D;
mem[16'hDC49] = 8'hA9;
mem[16'hDC4A] = 8'h2C;
mem[16'hDC4B] = 8'h18;
mem[16'hDC4C] = 8'h85;
mem[16'hDC4D] = 8'h0E;
mem[16'hDC4E] = 8'hA5;
mem[16'hDC4F] = 8'hB8;
mem[16'hDC50] = 8'hA4;
mem[16'hDC51] = 8'hB9;
mem[16'hDC52] = 8'h69;
mem[16'hDC53] = 8'h00;
mem[16'hDC54] = 8'h90;
mem[16'hDC55] = 8'h01;
mem[16'hDC56] = 8'hC8;
mem[16'hDC57] = 8'h20;
mem[16'hDC58] = 8'hED;
mem[16'hDC59] = 8'hE3;
mem[16'hDC5A] = 8'h20;
mem[16'hDC5B] = 8'h3D;
mem[16'hDC5C] = 8'hE7;
mem[16'hDC5D] = 8'h20;
mem[16'hDC5E] = 8'h7B;
mem[16'hDC5F] = 8'hDA;
mem[16'hDC60] = 8'h4C;
mem[16'hDC61] = 8'h72;
mem[16'hDC62] = 8'hDC;
mem[16'hDC63] = 8'h48;
mem[16'hDC64] = 8'hAD;
mem[16'hDC65] = 8'h00;
mem[16'hDC66] = 8'h02;
mem[16'hDC67] = 8'hF0;
mem[16'hDC68] = 8'h30;
mem[16'hDC69] = 8'h68;
mem[16'hDC6A] = 8'h20;
mem[16'hDC6B] = 8'h4A;
mem[16'hDC6C] = 8'hEC;
mem[16'hDC6D] = 8'hA5;
mem[16'hDC6E] = 8'h12;
mem[16'hDC6F] = 8'h20;
mem[16'hDC70] = 8'h63;
mem[16'hDC71] = 8'hDA;
mem[16'hDC72] = 8'h20;
mem[16'hDC73] = 8'hB7;
mem[16'hDC74] = 8'h00;
mem[16'hDC75] = 8'hF0;
mem[16'hDC76] = 8'h07;
mem[16'hDC77] = 8'hC9;
mem[16'hDC78] = 8'h2C;
mem[16'hDC79] = 8'hF0;
mem[16'hDC7A] = 8'h03;
mem[16'hDC7B] = 8'h4C;
mem[16'hDC7C] = 8'h71;
mem[16'hDC7D] = 8'hDB;
mem[16'hDC7E] = 8'hA5;
mem[16'hDC7F] = 8'hB8;
mem[16'hDC80] = 8'hA4;
mem[16'hDC81] = 8'hB9;
mem[16'hDC82] = 8'h85;
mem[16'hDC83] = 8'h7F;
mem[16'hDC84] = 8'h84;
mem[16'hDC85] = 8'h80;
mem[16'hDC86] = 8'hA5;
mem[16'hDC87] = 8'h87;
mem[16'hDC88] = 8'hA4;
mem[16'hDC89] = 8'h88;
mem[16'hDC8A] = 8'h85;
mem[16'hDC8B] = 8'hB8;
mem[16'hDC8C] = 8'h84;
mem[16'hDC8D] = 8'hB9;
mem[16'hDC8E] = 8'h20;
mem[16'hDC8F] = 8'hB7;
mem[16'hDC90] = 8'h00;
mem[16'hDC91] = 8'hF0;
mem[16'hDC92] = 8'h33;
mem[16'hDC93] = 8'h20;
mem[16'hDC94] = 8'hBE;
mem[16'hDC95] = 8'hDE;
mem[16'hDC96] = 8'h4C;
mem[16'hDC97] = 8'hF1;
mem[16'hDC98] = 8'hDB;
mem[16'hDC99] = 8'hA5;
mem[16'hDC9A] = 8'h15;
mem[16'hDC9B] = 8'hD0;
mem[16'hDC9C] = 8'hCC;
mem[16'hDC9D] = 8'h4C;
mem[16'hDC9E] = 8'h86;
mem[16'hDC9F] = 8'hDB;
mem[16'hDCA0] = 8'h20;
mem[16'hDCA1] = 8'hA3;
mem[16'hDCA2] = 8'hD9;
mem[16'hDCA3] = 8'hC8;
mem[16'hDCA4] = 8'hAA;
mem[16'hDCA5] = 8'hD0;
mem[16'hDCA6] = 8'h12;
mem[16'hDCA7] = 8'hA2;
mem[16'hDCA8] = 8'h2A;
mem[16'hDCA9] = 8'hC8;
mem[16'hDCAA] = 8'hB1;
mem[16'hDCAB] = 8'hB8;
mem[16'hDCAC] = 8'hF0;
mem[16'hDCAD] = 8'h5F;
mem[16'hDCAE] = 8'hC8;
mem[16'hDCAF] = 8'hB1;
mem[16'hDCB0] = 8'hB8;
mem[16'hDCB1] = 8'h85;
mem[16'hDCB2] = 8'h7B;
mem[16'hDCB3] = 8'hC8;
mem[16'hDCB4] = 8'hB1;
mem[16'hDCB5] = 8'hB8;
mem[16'hDCB6] = 8'hC8;
mem[16'hDCB7] = 8'h85;
mem[16'hDCB8] = 8'h7C;
mem[16'hDCB9] = 8'hB1;
mem[16'hDCBA] = 8'hB8;
mem[16'hDCBB] = 8'hAA;
mem[16'hDCBC] = 8'h20;
mem[16'hDCBD] = 8'h98;
mem[16'hDCBE] = 8'hD9;
mem[16'hDCBF] = 8'hE0;
mem[16'hDCC0] = 8'h83;
mem[16'hDCC1] = 8'hD0;
mem[16'hDCC2] = 8'hDD;
mem[16'hDCC3] = 8'h4C;
mem[16'hDCC4] = 8'h2B;
mem[16'hDCC5] = 8'hDC;
mem[16'hDCC6] = 8'hA5;
mem[16'hDCC7] = 8'h7F;
mem[16'hDCC8] = 8'hA4;
mem[16'hDCC9] = 8'h80;
mem[16'hDCCA] = 8'hA6;
mem[16'hDCCB] = 8'h15;
mem[16'hDCCC] = 8'h10;
mem[16'hDCCD] = 8'h03;
mem[16'hDCCE] = 8'h4C;
mem[16'hDCCF] = 8'h53;
mem[16'hDCD0] = 8'hD8;
mem[16'hDCD1] = 8'hA0;
mem[16'hDCD2] = 8'h00;
mem[16'hDCD3] = 8'hB1;
mem[16'hDCD4] = 8'h7F;
mem[16'hDCD5] = 8'hF0;
mem[16'hDCD6] = 8'h07;
mem[16'hDCD7] = 8'hA9;
mem[16'hDCD8] = 8'hDF;
mem[16'hDCD9] = 8'hA0;
mem[16'hDCDA] = 8'hDC;
mem[16'hDCDB] = 8'h4C;
mem[16'hDCDC] = 8'h3A;
mem[16'hDCDD] = 8'hDB;
mem[16'hDCDE] = 8'h60;
mem[16'hDCDF] = 8'h3F;
mem[16'hDCE0] = 8'h45;
mem[16'hDCE1] = 8'h58;
mem[16'hDCE2] = 8'h54;
mem[16'hDCE3] = 8'h52;
mem[16'hDCE4] = 8'h41;
mem[16'hDCE5] = 8'h20;
mem[16'hDCE6] = 8'h49;
mem[16'hDCE7] = 8'h47;
mem[16'hDCE8] = 8'h4E;
mem[16'hDCE9] = 8'h4F;
mem[16'hDCEA] = 8'h52;
mem[16'hDCEB] = 8'h45;
mem[16'hDCEC] = 8'h44;
mem[16'hDCED] = 8'h0D;
mem[16'hDCEE] = 8'h00;
mem[16'hDCEF] = 8'h3F;
mem[16'hDCF0] = 8'h52;
mem[16'hDCF1] = 8'h45;
mem[16'hDCF2] = 8'h45;
mem[16'hDCF3] = 8'h4E;
mem[16'hDCF4] = 8'h54;
mem[16'hDCF5] = 8'h45;
mem[16'hDCF6] = 8'h52;
mem[16'hDCF7] = 8'h0D;
mem[16'hDCF8] = 8'h00;
mem[16'hDCF9] = 8'hD0;
mem[16'hDCFA] = 8'h04;
mem[16'hDCFB] = 8'hA0;
mem[16'hDCFC] = 8'h00;
mem[16'hDCFD] = 8'hF0;
mem[16'hDCFE] = 8'h03;
mem[16'hDCFF] = 8'h20;
mem[16'hDD00] = 8'hE3;
mem[16'hDD01] = 8'hDF;
mem[16'hDD02] = 8'h85;
mem[16'hDD03] = 8'h85;
mem[16'hDD04] = 8'h84;
mem[16'hDD05] = 8'h86;
mem[16'hDD06] = 8'h20;
mem[16'hDD07] = 8'h65;
mem[16'hDD08] = 8'hD3;
mem[16'hDD09] = 8'hF0;
mem[16'hDD0A] = 8'h04;
mem[16'hDD0B] = 8'hA2;
mem[16'hDD0C] = 8'h00;
mem[16'hDD0D] = 8'hF0;
mem[16'hDD0E] = 8'h69;
mem[16'hDD0F] = 8'h9A;
mem[16'hDD10] = 8'hE8;
mem[16'hDD11] = 8'hE8;
mem[16'hDD12] = 8'hE8;
mem[16'hDD13] = 8'hE8;
mem[16'hDD14] = 8'h8A;
mem[16'hDD15] = 8'hE8;
mem[16'hDD16] = 8'hE8;
mem[16'hDD17] = 8'hE8;
mem[16'hDD18] = 8'hE8;
mem[16'hDD19] = 8'hE8;
mem[16'hDD1A] = 8'hE8;
mem[16'hDD1B] = 8'h86;
mem[16'hDD1C] = 8'h60;
mem[16'hDD1D] = 8'hA0;
mem[16'hDD1E] = 8'h01;
mem[16'hDD1F] = 8'h20;
mem[16'hDD20] = 8'hF9;
mem[16'hDD21] = 8'hEA;
mem[16'hDD22] = 8'hBA;
mem[16'hDD23] = 8'hBD;
mem[16'hDD24] = 8'h09;
mem[16'hDD25] = 8'h01;
mem[16'hDD26] = 8'h85;
mem[16'hDD27] = 8'hA2;
mem[16'hDD28] = 8'hA5;
mem[16'hDD29] = 8'h85;
mem[16'hDD2A] = 8'hA4;
mem[16'hDD2B] = 8'h86;
mem[16'hDD2C] = 8'h20;
mem[16'hDD2D] = 8'hBE;
mem[16'hDD2E] = 8'hE7;
mem[16'hDD2F] = 8'h20;
mem[16'hDD30] = 8'h27;
mem[16'hDD31] = 8'hEB;
mem[16'hDD32] = 8'hA0;
mem[16'hDD33] = 8'h01;
mem[16'hDD34] = 8'h20;
mem[16'hDD35] = 8'hB4;
mem[16'hDD36] = 8'hEB;
mem[16'hDD37] = 8'hBA;
mem[16'hDD38] = 8'h38;
mem[16'hDD39] = 8'hFD;
mem[16'hDD3A] = 8'h09;
mem[16'hDD3B] = 8'h01;
mem[16'hDD3C] = 8'hF0;
mem[16'hDD3D] = 8'h17;
mem[16'hDD3E] = 8'hBD;
mem[16'hDD3F] = 8'h0F;
mem[16'hDD40] = 8'h01;
mem[16'hDD41] = 8'h85;
mem[16'hDD42] = 8'h75;
mem[16'hDD43] = 8'hBD;
mem[16'hDD44] = 8'h10;
mem[16'hDD45] = 8'h01;
mem[16'hDD46] = 8'h85;
mem[16'hDD47] = 8'h76;
mem[16'hDD48] = 8'hBD;
mem[16'hDD49] = 8'h12;
mem[16'hDD4A] = 8'h01;
mem[16'hDD4B] = 8'h85;
mem[16'hDD4C] = 8'hB8;
mem[16'hDD4D] = 8'hBD;
mem[16'hDD4E] = 8'h11;
mem[16'hDD4F] = 8'h01;
mem[16'hDD50] = 8'h85;
mem[16'hDD51] = 8'hB9;
mem[16'hDD52] = 8'h4C;
mem[16'hDD53] = 8'hD2;
mem[16'hDD54] = 8'hD7;
mem[16'hDD55] = 8'h8A;
mem[16'hDD56] = 8'h69;
mem[16'hDD57] = 8'h11;
mem[16'hDD58] = 8'hAA;
mem[16'hDD59] = 8'h9A;
mem[16'hDD5A] = 8'h20;
mem[16'hDD5B] = 8'hB7;
mem[16'hDD5C] = 8'h00;
mem[16'hDD5D] = 8'hC9;
mem[16'hDD5E] = 8'h2C;
mem[16'hDD5F] = 8'hD0;
mem[16'hDD60] = 8'hF1;
mem[16'hDD61] = 8'h20;
mem[16'hDD62] = 8'hB1;
mem[16'hDD63] = 8'h00;
mem[16'hDD64] = 8'h20;
mem[16'hDD65] = 8'hFF;
mem[16'hDD66] = 8'hDC;
mem[16'hDD67] = 8'h20;
mem[16'hDD68] = 8'h7B;
mem[16'hDD69] = 8'hDD;
mem[16'hDD6A] = 8'h18;
mem[16'hDD6B] = 8'h24;
mem[16'hDD6C] = 8'h38;
mem[16'hDD6D] = 8'h24;
mem[16'hDD6E] = 8'h11;
mem[16'hDD6F] = 8'h30;
mem[16'hDD70] = 8'h03;
mem[16'hDD71] = 8'hB0;
mem[16'hDD72] = 8'h03;
mem[16'hDD73] = 8'h60;
mem[16'hDD74] = 8'hB0;
mem[16'hDD75] = 8'hFD;
mem[16'hDD76] = 8'hA2;
mem[16'hDD77] = 8'hA3;
mem[16'hDD78] = 8'h4C;
mem[16'hDD79] = 8'h12;
mem[16'hDD7A] = 8'hD4;
mem[16'hDD7B] = 8'hA6;
mem[16'hDD7C] = 8'hB8;
mem[16'hDD7D] = 8'hD0;
mem[16'hDD7E] = 8'h02;
mem[16'hDD7F] = 8'hC6;
mem[16'hDD80] = 8'hB9;
mem[16'hDD81] = 8'hC6;
mem[16'hDD82] = 8'hB8;
mem[16'hDD83] = 8'hA2;
mem[16'hDD84] = 8'h00;
mem[16'hDD85] = 8'h24;
mem[16'hDD86] = 8'h48;
mem[16'hDD87] = 8'h8A;
mem[16'hDD88] = 8'h48;
mem[16'hDD89] = 8'hA9;
mem[16'hDD8A] = 8'h01;
mem[16'hDD8B] = 8'h20;
mem[16'hDD8C] = 8'hD6;
mem[16'hDD8D] = 8'hD3;
mem[16'hDD8E] = 8'h20;
mem[16'hDD8F] = 8'h60;
mem[16'hDD90] = 8'hDE;
mem[16'hDD91] = 8'hA9;
mem[16'hDD92] = 8'h00;
mem[16'hDD93] = 8'h85;
mem[16'hDD94] = 8'h89;
mem[16'hDD95] = 8'h20;
mem[16'hDD96] = 8'hB7;
mem[16'hDD97] = 8'h00;
mem[16'hDD98] = 8'h38;
mem[16'hDD99] = 8'hE9;
mem[16'hDD9A] = 8'hCF;
mem[16'hDD9B] = 8'h90;
mem[16'hDD9C] = 8'h17;
mem[16'hDD9D] = 8'hC9;
mem[16'hDD9E] = 8'h03;
mem[16'hDD9F] = 8'hB0;
mem[16'hDDA0] = 8'h13;
mem[16'hDDA1] = 8'hC9;
mem[16'hDDA2] = 8'h01;
mem[16'hDDA3] = 8'h2A;
mem[16'hDDA4] = 8'h49;
mem[16'hDDA5] = 8'h01;
mem[16'hDDA6] = 8'h45;
mem[16'hDDA7] = 8'h89;
mem[16'hDDA8] = 8'hC5;
mem[16'hDDA9] = 8'h89;
mem[16'hDDAA] = 8'h90;
mem[16'hDDAB] = 8'h61;
mem[16'hDDAC] = 8'h85;
mem[16'hDDAD] = 8'h89;
mem[16'hDDAE] = 8'h20;
mem[16'hDDAF] = 8'hB1;
mem[16'hDDB0] = 8'h00;
mem[16'hDDB1] = 8'h4C;
mem[16'hDDB2] = 8'h98;
mem[16'hDDB3] = 8'hDD;
mem[16'hDDB4] = 8'hA6;
mem[16'hDDB5] = 8'h89;
mem[16'hDDB6] = 8'hD0;
mem[16'hDDB7] = 8'h2C;
mem[16'hDDB8] = 8'hB0;
mem[16'hDDB9] = 8'h7B;
mem[16'hDDBA] = 8'h69;
mem[16'hDDBB] = 8'h07;
mem[16'hDDBC] = 8'h90;
mem[16'hDDBD] = 8'h77;
mem[16'hDDBE] = 8'h65;
mem[16'hDDBF] = 8'h11;
mem[16'hDDC0] = 8'hD0;
mem[16'hDDC1] = 8'h03;
mem[16'hDDC2] = 8'h4C;
mem[16'hDDC3] = 8'h97;
mem[16'hDDC4] = 8'hE5;
mem[16'hDDC5] = 8'h69;
mem[16'hDDC6] = 8'hFF;
mem[16'hDDC7] = 8'h85;
mem[16'hDDC8] = 8'h5E;
mem[16'hDDC9] = 8'h0A;
mem[16'hDDCA] = 8'h65;
mem[16'hDDCB] = 8'h5E;
mem[16'hDDCC] = 8'hA8;
mem[16'hDDCD] = 8'h68;
mem[16'hDDCE] = 8'hD9;
mem[16'hDDCF] = 8'hB2;
mem[16'hDDD0] = 8'hD0;
mem[16'hDDD1] = 8'hB0;
mem[16'hDDD2] = 8'h67;
mem[16'hDDD3] = 8'h20;
mem[16'hDDD4] = 8'h6A;
mem[16'hDDD5] = 8'hDD;
mem[16'hDDD6] = 8'h48;
mem[16'hDDD7] = 8'h20;
mem[16'hDDD8] = 8'hFD;
mem[16'hDDD9] = 8'hDD;
mem[16'hDDDA] = 8'h68;
mem[16'hDDDB] = 8'hA4;
mem[16'hDDDC] = 8'h87;
mem[16'hDDDD] = 8'h10;
mem[16'hDDDE] = 8'h17;
mem[16'hDDDF] = 8'hAA;
mem[16'hDDE0] = 8'hF0;
mem[16'hDDE1] = 8'h56;
mem[16'hDDE2] = 8'hD0;
mem[16'hDDE3] = 8'h5F;
mem[16'hDDE4] = 8'h46;
mem[16'hDDE5] = 8'h11;
mem[16'hDDE6] = 8'h8A;
mem[16'hDDE7] = 8'h2A;
mem[16'hDDE8] = 8'hA6;
mem[16'hDDE9] = 8'hB8;
mem[16'hDDEA] = 8'hD0;
mem[16'hDDEB] = 8'h02;
mem[16'hDDEC] = 8'hC6;
mem[16'hDDED] = 8'hB9;
mem[16'hDDEE] = 8'hC6;
mem[16'hDDEF] = 8'hB8;
mem[16'hDDF0] = 8'hA0;
mem[16'hDDF1] = 8'h1B;
mem[16'hDDF2] = 8'h85;
mem[16'hDDF3] = 8'h89;
mem[16'hDDF4] = 8'hD0;
mem[16'hDDF5] = 8'hD7;
mem[16'hDDF6] = 8'hD9;
mem[16'hDDF7] = 8'hB2;
mem[16'hDDF8] = 8'hD0;
mem[16'hDDF9] = 8'hB0;
mem[16'hDDFA] = 8'h48;
mem[16'hDDFB] = 8'h90;
mem[16'hDDFC] = 8'hD9;
mem[16'hDDFD] = 8'hB9;
mem[16'hDDFE] = 8'hB4;
mem[16'hDDFF] = 8'hD0;
mem[16'hDE00] = 8'h48;
mem[16'hDE01] = 8'hB9;
mem[16'hDE02] = 8'hB3;
mem[16'hDE03] = 8'hD0;
mem[16'hDE04] = 8'h48;
mem[16'hDE05] = 8'h20;
mem[16'hDE06] = 8'h10;
mem[16'hDE07] = 8'hDE;
mem[16'hDE08] = 8'hA5;
mem[16'hDE09] = 8'h89;
mem[16'hDE0A] = 8'h4C;
mem[16'hDE0B] = 8'h86;
mem[16'hDE0C] = 8'hDD;
mem[16'hDE0D] = 8'h4C;
mem[16'hDE0E] = 8'hC9;
mem[16'hDE0F] = 8'hDE;
mem[16'hDE10] = 8'hA5;
mem[16'hDE11] = 8'hA2;
mem[16'hDE12] = 8'hBE;
mem[16'hDE13] = 8'hB2;
mem[16'hDE14] = 8'hD0;
mem[16'hDE15] = 8'hA8;
mem[16'hDE16] = 8'h68;
mem[16'hDE17] = 8'h85;
mem[16'hDE18] = 8'h5E;
mem[16'hDE19] = 8'hE6;
mem[16'hDE1A] = 8'h5E;
mem[16'hDE1B] = 8'h68;
mem[16'hDE1C] = 8'h85;
mem[16'hDE1D] = 8'h5F;
mem[16'hDE1E] = 8'h98;
mem[16'hDE1F] = 8'h48;
mem[16'hDE20] = 8'h20;
mem[16'hDE21] = 8'h72;
mem[16'hDE22] = 8'hEB;
mem[16'hDE23] = 8'hA5;
mem[16'hDE24] = 8'hA1;
mem[16'hDE25] = 8'h48;
mem[16'hDE26] = 8'hA5;
mem[16'hDE27] = 8'hA0;
mem[16'hDE28] = 8'h48;
mem[16'hDE29] = 8'hA5;
mem[16'hDE2A] = 8'h9F;
mem[16'hDE2B] = 8'h48;
mem[16'hDE2C] = 8'hA5;
mem[16'hDE2D] = 8'h9E;
mem[16'hDE2E] = 8'h48;
mem[16'hDE2F] = 8'hA5;
mem[16'hDE30] = 8'h9D;
mem[16'hDE31] = 8'h48;
mem[16'hDE32] = 8'h6C;
mem[16'hDE33] = 8'h5E;
mem[16'hDE34] = 8'h00;
mem[16'hDE35] = 8'hA0;
mem[16'hDE36] = 8'hFF;
mem[16'hDE37] = 8'h68;
mem[16'hDE38] = 8'hF0;
mem[16'hDE39] = 8'h23;
mem[16'hDE3A] = 8'hC9;
mem[16'hDE3B] = 8'h64;
mem[16'hDE3C] = 8'hF0;
mem[16'hDE3D] = 8'h03;
mem[16'hDE3E] = 8'h20;
mem[16'hDE3F] = 8'h6A;
mem[16'hDE40] = 8'hDD;
mem[16'hDE41] = 8'h84;
mem[16'hDE42] = 8'h87;
mem[16'hDE43] = 8'h68;
mem[16'hDE44] = 8'h4A;
mem[16'hDE45] = 8'h85;
mem[16'hDE46] = 8'h16;
mem[16'hDE47] = 8'h68;
mem[16'hDE48] = 8'h85;
mem[16'hDE49] = 8'hA5;
mem[16'hDE4A] = 8'h68;
mem[16'hDE4B] = 8'h85;
mem[16'hDE4C] = 8'hA6;
mem[16'hDE4D] = 8'h68;
mem[16'hDE4E] = 8'h85;
mem[16'hDE4F] = 8'hA7;
mem[16'hDE50] = 8'h68;
mem[16'hDE51] = 8'h85;
mem[16'hDE52] = 8'hA8;
mem[16'hDE53] = 8'h68;
mem[16'hDE54] = 8'h85;
mem[16'hDE55] = 8'hA9;
mem[16'hDE56] = 8'h68;
mem[16'hDE57] = 8'h85;
mem[16'hDE58] = 8'hAA;
mem[16'hDE59] = 8'h45;
mem[16'hDE5A] = 8'hA2;
mem[16'hDE5B] = 8'h85;
mem[16'hDE5C] = 8'hAB;
mem[16'hDE5D] = 8'hA5;
mem[16'hDE5E] = 8'h9D;
mem[16'hDE5F] = 8'h60;
mem[16'hDE60] = 8'hA9;
mem[16'hDE61] = 8'h00;
mem[16'hDE62] = 8'h85;
mem[16'hDE63] = 8'h11;
mem[16'hDE64] = 8'h20;
mem[16'hDE65] = 8'hB1;
mem[16'hDE66] = 8'h00;
mem[16'hDE67] = 8'hB0;
mem[16'hDE68] = 8'h03;
mem[16'hDE69] = 8'h4C;
mem[16'hDE6A] = 8'h4A;
mem[16'hDE6B] = 8'hEC;
mem[16'hDE6C] = 8'h20;
mem[16'hDE6D] = 8'h7D;
mem[16'hDE6E] = 8'hE0;
mem[16'hDE6F] = 8'hB0;
mem[16'hDE70] = 8'h64;
mem[16'hDE71] = 8'hC9;
mem[16'hDE72] = 8'h2E;
mem[16'hDE73] = 8'hF0;
mem[16'hDE74] = 8'hF4;
mem[16'hDE75] = 8'hC9;
mem[16'hDE76] = 8'hC9;
mem[16'hDE77] = 8'hF0;
mem[16'hDE78] = 8'h55;
mem[16'hDE79] = 8'hC9;
mem[16'hDE7A] = 8'hC8;
mem[16'hDE7B] = 8'hF0;
mem[16'hDE7C] = 8'hE7;
mem[16'hDE7D] = 8'hC9;
mem[16'hDE7E] = 8'h22;
mem[16'hDE7F] = 8'hD0;
mem[16'hDE80] = 8'h0F;
mem[16'hDE81] = 8'hA5;
mem[16'hDE82] = 8'hB8;
mem[16'hDE83] = 8'hA4;
mem[16'hDE84] = 8'hB9;
mem[16'hDE85] = 8'h69;
mem[16'hDE86] = 8'h00;
mem[16'hDE87] = 8'h90;
mem[16'hDE88] = 8'h01;
mem[16'hDE89] = 8'hC8;
mem[16'hDE8A] = 8'h20;
mem[16'hDE8B] = 8'hE7;
mem[16'hDE8C] = 8'hE3;
mem[16'hDE8D] = 8'h4C;
mem[16'hDE8E] = 8'h3D;
mem[16'hDE8F] = 8'hE7;
mem[16'hDE90] = 8'hC9;
mem[16'hDE91] = 8'hC6;
mem[16'hDE92] = 8'hD0;
mem[16'hDE93] = 8'h10;
mem[16'hDE94] = 8'hA0;
mem[16'hDE95] = 8'h18;
mem[16'hDE96] = 8'hD0;
mem[16'hDE97] = 8'h38;
mem[16'hDE98] = 8'hA5;
mem[16'hDE99] = 8'h9D;
mem[16'hDE9A] = 8'hD0;
mem[16'hDE9B] = 8'h03;
mem[16'hDE9C] = 8'hA0;
mem[16'hDE9D] = 8'h01;
mem[16'hDE9E] = 8'h2C;
mem[16'hDE9F] = 8'hA0;
mem[16'hDEA0] = 8'h00;
mem[16'hDEA1] = 8'h4C;
mem[16'hDEA2] = 8'h01;
mem[16'hDEA3] = 8'hE3;
mem[16'hDEA4] = 8'hC9;
mem[16'hDEA5] = 8'hC2;
mem[16'hDEA6] = 8'hD0;
mem[16'hDEA7] = 8'h03;
mem[16'hDEA8] = 8'h4C;
mem[16'hDEA9] = 8'h54;
mem[16'hDEAA] = 8'hE3;
mem[16'hDEAB] = 8'hC9;
mem[16'hDEAC] = 8'hD2;
mem[16'hDEAD] = 8'h90;
mem[16'hDEAE] = 8'h03;
mem[16'hDEAF] = 8'h4C;
mem[16'hDEB0] = 8'h0C;
mem[16'hDEB1] = 8'hDF;
mem[16'hDEB2] = 8'h20;
mem[16'hDEB3] = 8'hBB;
mem[16'hDEB4] = 8'hDE;
mem[16'hDEB5] = 8'h20;
mem[16'hDEB6] = 8'h7B;
mem[16'hDEB7] = 8'hDD;
mem[16'hDEB8] = 8'hA9;
mem[16'hDEB9] = 8'h29;
mem[16'hDEBA] = 8'h2C;
mem[16'hDEBB] = 8'hA9;
mem[16'hDEBC] = 8'h28;
mem[16'hDEBD] = 8'h2C;
mem[16'hDEBE] = 8'hA9;
mem[16'hDEBF] = 8'h2C;
mem[16'hDEC0] = 8'hA0;
mem[16'hDEC1] = 8'h00;
mem[16'hDEC2] = 8'hD1;
mem[16'hDEC3] = 8'hB8;
mem[16'hDEC4] = 8'hD0;
mem[16'hDEC5] = 8'h03;
mem[16'hDEC6] = 8'h4C;
mem[16'hDEC7] = 8'hB1;
mem[16'hDEC8] = 8'h00;
mem[16'hDEC9] = 8'hA2;
mem[16'hDECA] = 8'h10;
mem[16'hDECB] = 8'h4C;
mem[16'hDECC] = 8'h12;
mem[16'hDECD] = 8'hD4;
mem[16'hDECE] = 8'hA0;
mem[16'hDECF] = 8'h15;
mem[16'hDED0] = 8'h68;
mem[16'hDED1] = 8'h68;
mem[16'hDED2] = 8'h4C;
mem[16'hDED3] = 8'hD7;
mem[16'hDED4] = 8'hDD;
mem[16'hDED5] = 8'h20;
mem[16'hDED6] = 8'hE3;
mem[16'hDED7] = 8'hDF;
mem[16'hDED8] = 8'h85;
mem[16'hDED9] = 8'hA0;
mem[16'hDEDA] = 8'h84;
mem[16'hDEDB] = 8'hA1;
mem[16'hDEDC] = 8'hA6;
mem[16'hDEDD] = 8'h11;
mem[16'hDEDE] = 8'hF0;
mem[16'hDEDF] = 8'h05;
mem[16'hDEE0] = 8'hA2;
mem[16'hDEE1] = 8'h00;
mem[16'hDEE2] = 8'h86;
mem[16'hDEE3] = 8'hAC;
mem[16'hDEE4] = 8'h60;
mem[16'hDEE5] = 8'hA6;
mem[16'hDEE6] = 8'h12;
mem[16'hDEE7] = 8'h10;
mem[16'hDEE8] = 8'h0D;
mem[16'hDEE9] = 8'hA0;
mem[16'hDEEA] = 8'h00;
mem[16'hDEEB] = 8'hB1;
mem[16'hDEEC] = 8'hA0;
mem[16'hDEED] = 8'hAA;
mem[16'hDEEE] = 8'hC8;
mem[16'hDEEF] = 8'hB1;
mem[16'hDEF0] = 8'hA0;
mem[16'hDEF1] = 8'hA8;
mem[16'hDEF2] = 8'h8A;
mem[16'hDEF3] = 8'h4C;
mem[16'hDEF4] = 8'hF2;
mem[16'hDEF5] = 8'hE2;
mem[16'hDEF6] = 8'h4C;
mem[16'hDEF7] = 8'hF9;
mem[16'hDEF8] = 8'hEA;
mem[16'hDEF9] = 8'h20;
mem[16'hDEFA] = 8'hB1;
mem[16'hDEFB] = 8'h00;
mem[16'hDEFC] = 8'h20;
mem[16'hDEFD] = 8'hEC;
mem[16'hDEFE] = 8'hF1;
mem[16'hDEFF] = 8'h8A;
mem[16'hDF00] = 8'hA4;
mem[16'hDF01] = 8'hF0;
mem[16'hDF02] = 8'h20;
mem[16'hDF03] = 8'h71;
mem[16'hDF04] = 8'hF8;
mem[16'hDF05] = 8'hA8;
mem[16'hDF06] = 8'h20;
mem[16'hDF07] = 8'h01;
mem[16'hDF08] = 8'hE3;
mem[16'hDF09] = 8'h4C;
mem[16'hDF0A] = 8'hB8;
mem[16'hDF0B] = 8'hDE;
mem[16'hDF0C] = 8'hC9;
mem[16'hDF0D] = 8'hD7;
mem[16'hDF0E] = 8'hF0;
mem[16'hDF0F] = 8'hE9;
mem[16'hDF10] = 8'h0A;
mem[16'hDF11] = 8'h48;
mem[16'hDF12] = 8'hAA;
mem[16'hDF13] = 8'h20;
mem[16'hDF14] = 8'hB1;
mem[16'hDF15] = 8'h00;
mem[16'hDF16] = 8'hE0;
mem[16'hDF17] = 8'hCF;
mem[16'hDF18] = 8'h90;
mem[16'hDF19] = 8'h20;
mem[16'hDF1A] = 8'h20;
mem[16'hDF1B] = 8'hBB;
mem[16'hDF1C] = 8'hDE;
mem[16'hDF1D] = 8'h20;
mem[16'hDF1E] = 8'h7B;
mem[16'hDF1F] = 8'hDD;
mem[16'hDF20] = 8'h20;
mem[16'hDF21] = 8'hBE;
mem[16'hDF22] = 8'hDE;
mem[16'hDF23] = 8'h20;
mem[16'hDF24] = 8'h6C;
mem[16'hDF25] = 8'hDD;
mem[16'hDF26] = 8'h68;
mem[16'hDF27] = 8'hAA;
mem[16'hDF28] = 8'hA5;
mem[16'hDF29] = 8'hA1;
mem[16'hDF2A] = 8'h48;
mem[16'hDF2B] = 8'hA5;
mem[16'hDF2C] = 8'hA0;
mem[16'hDF2D] = 8'h48;
mem[16'hDF2E] = 8'h8A;
mem[16'hDF2F] = 8'h48;
mem[16'hDF30] = 8'h20;
mem[16'hDF31] = 8'hF8;
mem[16'hDF32] = 8'hE6;
mem[16'hDF33] = 8'h68;
mem[16'hDF34] = 8'hA8;
mem[16'hDF35] = 8'h8A;
mem[16'hDF36] = 8'h48;
mem[16'hDF37] = 8'h4C;
mem[16'hDF38] = 8'h3F;
mem[16'hDF39] = 8'hDF;
mem[16'hDF3A] = 8'h20;
mem[16'hDF3B] = 8'hB2;
mem[16'hDF3C] = 8'hDE;
mem[16'hDF3D] = 8'h68;
mem[16'hDF3E] = 8'hA8;
mem[16'hDF3F] = 8'hB9;
mem[16'hDF40] = 8'hDC;
mem[16'hDF41] = 8'hCF;
mem[16'hDF42] = 8'h85;
mem[16'hDF43] = 8'h91;
mem[16'hDF44] = 8'hB9;
mem[16'hDF45] = 8'hDD;
mem[16'hDF46] = 8'hCF;
mem[16'hDF47] = 8'h85;
mem[16'hDF48] = 8'h92;
mem[16'hDF49] = 8'h20;
mem[16'hDF4A] = 8'h90;
mem[16'hDF4B] = 8'h00;
mem[16'hDF4C] = 8'h4C;
mem[16'hDF4D] = 8'h6A;
mem[16'hDF4E] = 8'hDD;
mem[16'hDF4F] = 8'hA5;
mem[16'hDF50] = 8'hA5;
mem[16'hDF51] = 8'h05;
mem[16'hDF52] = 8'h9D;
mem[16'hDF53] = 8'hD0;
mem[16'hDF54] = 8'h0B;
mem[16'hDF55] = 8'hA5;
mem[16'hDF56] = 8'hA5;
mem[16'hDF57] = 8'hF0;
mem[16'hDF58] = 8'h04;
mem[16'hDF59] = 8'hA5;
mem[16'hDF5A] = 8'h9D;
mem[16'hDF5B] = 8'hD0;
mem[16'hDF5C] = 8'h03;
mem[16'hDF5D] = 8'hA0;
mem[16'hDF5E] = 8'h00;
mem[16'hDF5F] = 8'h2C;
mem[16'hDF60] = 8'hA0;
mem[16'hDF61] = 8'h01;
mem[16'hDF62] = 8'h4C;
mem[16'hDF63] = 8'h01;
mem[16'hDF64] = 8'hE3;
mem[16'hDF65] = 8'h20;
mem[16'hDF66] = 8'h6D;
mem[16'hDF67] = 8'hDD;
mem[16'hDF68] = 8'hB0;
mem[16'hDF69] = 8'h13;
mem[16'hDF6A] = 8'hA5;
mem[16'hDF6B] = 8'hAA;
mem[16'hDF6C] = 8'h09;
mem[16'hDF6D] = 8'h7F;
mem[16'hDF6E] = 8'h25;
mem[16'hDF6F] = 8'hA6;
mem[16'hDF70] = 8'h85;
mem[16'hDF71] = 8'hA6;
mem[16'hDF72] = 8'hA9;
mem[16'hDF73] = 8'hA5;
mem[16'hDF74] = 8'hA0;
mem[16'hDF75] = 8'h00;
mem[16'hDF76] = 8'h20;
mem[16'hDF77] = 8'hB2;
mem[16'hDF78] = 8'hEB;
mem[16'hDF79] = 8'hAA;
mem[16'hDF7A] = 8'h4C;
mem[16'hDF7B] = 8'hB0;
mem[16'hDF7C] = 8'hDF;
mem[16'hDF7D] = 8'hA9;
mem[16'hDF7E] = 8'h00;
mem[16'hDF7F] = 8'h85;
mem[16'hDF80] = 8'h11;
mem[16'hDF81] = 8'hC6;
mem[16'hDF82] = 8'h89;
mem[16'hDF83] = 8'h20;
mem[16'hDF84] = 8'h00;
mem[16'hDF85] = 8'hE6;
mem[16'hDF86] = 8'h85;
mem[16'hDF87] = 8'h9D;
mem[16'hDF88] = 8'h86;
mem[16'hDF89] = 8'h9E;
mem[16'hDF8A] = 8'h84;
mem[16'hDF8B] = 8'h9F;
mem[16'hDF8C] = 8'hA5;
mem[16'hDF8D] = 8'hA8;
mem[16'hDF8E] = 8'hA4;
mem[16'hDF8F] = 8'hA9;
mem[16'hDF90] = 8'h20;
mem[16'hDF91] = 8'h04;
mem[16'hDF92] = 8'hE6;
mem[16'hDF93] = 8'h86;
mem[16'hDF94] = 8'hA8;
mem[16'hDF95] = 8'h84;
mem[16'hDF96] = 8'hA9;
mem[16'hDF97] = 8'hAA;
mem[16'hDF98] = 8'h38;
mem[16'hDF99] = 8'hE5;
mem[16'hDF9A] = 8'h9D;
mem[16'hDF9B] = 8'hF0;
mem[16'hDF9C] = 8'h08;
mem[16'hDF9D] = 8'hA9;
mem[16'hDF9E] = 8'h01;
mem[16'hDF9F] = 8'h90;
mem[16'hDFA0] = 8'h04;
mem[16'hDFA1] = 8'hA6;
mem[16'hDFA2] = 8'h9D;
mem[16'hDFA3] = 8'hA9;
mem[16'hDFA4] = 8'hFF;
mem[16'hDFA5] = 8'h85;
mem[16'hDFA6] = 8'hA2;
mem[16'hDFA7] = 8'hA0;
mem[16'hDFA8] = 8'hFF;
mem[16'hDFA9] = 8'hE8;
mem[16'hDFAA] = 8'hC8;
mem[16'hDFAB] = 8'hCA;
mem[16'hDFAC] = 8'hD0;
mem[16'hDFAD] = 8'h07;
mem[16'hDFAE] = 8'hA6;
mem[16'hDFAF] = 8'hA2;
mem[16'hDFB0] = 8'h30;
mem[16'hDFB1] = 8'h0F;
mem[16'hDFB2] = 8'h18;
mem[16'hDFB3] = 8'h90;
mem[16'hDFB4] = 8'h0C;
mem[16'hDFB5] = 8'hB1;
mem[16'hDFB6] = 8'hA8;
mem[16'hDFB7] = 8'hD1;
mem[16'hDFB8] = 8'h9E;
mem[16'hDFB9] = 8'hF0;
mem[16'hDFBA] = 8'hEF;
mem[16'hDFBB] = 8'hA2;
mem[16'hDFBC] = 8'hFF;
mem[16'hDFBD] = 8'hB0;
mem[16'hDFBE] = 8'h02;
mem[16'hDFBF] = 8'hA2;
mem[16'hDFC0] = 8'h01;
mem[16'hDFC1] = 8'hE8;
mem[16'hDFC2] = 8'h8A;
mem[16'hDFC3] = 8'h2A;
mem[16'hDFC4] = 8'h25;
mem[16'hDFC5] = 8'h16;
mem[16'hDFC6] = 8'hF0;
mem[16'hDFC7] = 8'h02;
mem[16'hDFC8] = 8'hA9;
mem[16'hDFC9] = 8'h01;
mem[16'hDFCA] = 8'h4C;
mem[16'hDFCB] = 8'h93;
mem[16'hDFCC] = 8'hEB;
mem[16'hDFCD] = 8'h20;
mem[16'hDFCE] = 8'hFB;
mem[16'hDFCF] = 8'hE6;
mem[16'hDFD0] = 8'h20;
mem[16'hDFD1] = 8'h1E;
mem[16'hDFD2] = 8'hFB;
mem[16'hDFD3] = 8'h4C;
mem[16'hDFD4] = 8'h01;
mem[16'hDFD5] = 8'hE3;
mem[16'hDFD6] = 8'h20;
mem[16'hDFD7] = 8'hBE;
mem[16'hDFD8] = 8'hDE;
mem[16'hDFD9] = 8'hAA;
mem[16'hDFDA] = 8'h20;
mem[16'hDFDB] = 8'hE8;
mem[16'hDFDC] = 8'hDF;
mem[16'hDFDD] = 8'h20;
mem[16'hDFDE] = 8'hB7;
mem[16'hDFDF] = 8'h00;
mem[16'hDFE0] = 8'hD0;
mem[16'hDFE1] = 8'hF4;
mem[16'hDFE2] = 8'h60;
mem[16'hDFE3] = 8'hA2;
mem[16'hDFE4] = 8'h00;
mem[16'hDFE5] = 8'h20;
mem[16'hDFE6] = 8'hB7;
mem[16'hDFE7] = 8'h00;
mem[16'hDFE8] = 8'h86;
mem[16'hDFE9] = 8'h10;
mem[16'hDFEA] = 8'h85;
mem[16'hDFEB] = 8'h81;
mem[16'hDFEC] = 8'h20;
mem[16'hDFED] = 8'hB7;
mem[16'hDFEE] = 8'h00;
mem[16'hDFEF] = 8'h20;
mem[16'hDFF0] = 8'h7D;
mem[16'hDFF1] = 8'hE0;
mem[16'hDFF2] = 8'hB0;
mem[16'hDFF3] = 8'h03;
mem[16'hDFF4] = 8'h4C;
mem[16'hDFF5] = 8'hC9;
mem[16'hDFF6] = 8'hDE;
mem[16'hDFF7] = 8'hA2;
mem[16'hDFF8] = 8'h00;
mem[16'hDFF9] = 8'h86;
mem[16'hDFFA] = 8'h11;
mem[16'hDFFB] = 8'h86;
mem[16'hDFFC] = 8'h12;
mem[16'hDFFD] = 8'h4C;
mem[16'hDFFE] = 8'h07;
mem[16'hDFFF] = 8'hE0;
mem[16'hE000] = 8'h4C;
mem[16'hE001] = 8'h28;
mem[16'hE002] = 8'hF1;
mem[16'hE003] = 8'h4C;
mem[16'hE004] = 8'h3C;
mem[16'hE005] = 8'hD4;
mem[16'hE006] = 8'h00;
mem[16'hE007] = 8'h20;
mem[16'hE008] = 8'hB1;
mem[16'hE009] = 8'h00;
mem[16'hE00A] = 8'h90;
mem[16'hE00B] = 8'h05;
mem[16'hE00C] = 8'h20;
mem[16'hE00D] = 8'h7D;
mem[16'hE00E] = 8'hE0;
mem[16'hE00F] = 8'h90;
mem[16'hE010] = 8'h0B;
mem[16'hE011] = 8'hAA;
mem[16'hE012] = 8'h20;
mem[16'hE013] = 8'hB1;
mem[16'hE014] = 8'h00;
mem[16'hE015] = 8'h90;
mem[16'hE016] = 8'hFB;
mem[16'hE017] = 8'h20;
mem[16'hE018] = 8'h7D;
mem[16'hE019] = 8'hE0;
mem[16'hE01A] = 8'hB0;
mem[16'hE01B] = 8'hF6;
mem[16'hE01C] = 8'hC9;
mem[16'hE01D] = 8'h24;
mem[16'hE01E] = 8'hD0;
mem[16'hE01F] = 8'h06;
mem[16'hE020] = 8'hA9;
mem[16'hE021] = 8'hFF;
mem[16'hE022] = 8'h85;
mem[16'hE023] = 8'h11;
mem[16'hE024] = 8'hD0;
mem[16'hE025] = 8'h10;
mem[16'hE026] = 8'hC9;
mem[16'hE027] = 8'h25;
mem[16'hE028] = 8'hD0;
mem[16'hE029] = 8'h13;
mem[16'hE02A] = 8'hA5;
mem[16'hE02B] = 8'h14;
mem[16'hE02C] = 8'h30;
mem[16'hE02D] = 8'hC6;
mem[16'hE02E] = 8'hA9;
mem[16'hE02F] = 8'h80;
mem[16'hE030] = 8'h85;
mem[16'hE031] = 8'h12;
mem[16'hE032] = 8'h05;
mem[16'hE033] = 8'h81;
mem[16'hE034] = 8'h85;
mem[16'hE035] = 8'h81;
mem[16'hE036] = 8'h8A;
mem[16'hE037] = 8'h09;
mem[16'hE038] = 8'h80;
mem[16'hE039] = 8'hAA;
mem[16'hE03A] = 8'h20;
mem[16'hE03B] = 8'hB1;
mem[16'hE03C] = 8'h00;
mem[16'hE03D] = 8'h86;
mem[16'hE03E] = 8'h82;
mem[16'hE03F] = 8'h38;
mem[16'hE040] = 8'h05;
mem[16'hE041] = 8'h14;
mem[16'hE042] = 8'hE9;
mem[16'hE043] = 8'h28;
mem[16'hE044] = 8'hD0;
mem[16'hE045] = 8'h03;
mem[16'hE046] = 8'h4C;
mem[16'hE047] = 8'h1E;
mem[16'hE048] = 8'hE1;
mem[16'hE049] = 8'h24;
mem[16'hE04A] = 8'h14;
mem[16'hE04B] = 8'h30;
mem[16'hE04C] = 8'h02;
mem[16'hE04D] = 8'h70;
mem[16'hE04E] = 8'hF7;
mem[16'hE04F] = 8'hA9;
mem[16'hE050] = 8'h00;
mem[16'hE051] = 8'h85;
mem[16'hE052] = 8'h14;
mem[16'hE053] = 8'hA5;
mem[16'hE054] = 8'h69;
mem[16'hE055] = 8'hA6;
mem[16'hE056] = 8'h6A;
mem[16'hE057] = 8'hA0;
mem[16'hE058] = 8'h00;
mem[16'hE059] = 8'h86;
mem[16'hE05A] = 8'h9C;
mem[16'hE05B] = 8'h85;
mem[16'hE05C] = 8'h9B;
mem[16'hE05D] = 8'hE4;
mem[16'hE05E] = 8'h6C;
mem[16'hE05F] = 8'hD0;
mem[16'hE060] = 8'h04;
mem[16'hE061] = 8'hC5;
mem[16'hE062] = 8'h6B;
mem[16'hE063] = 8'hF0;
mem[16'hE064] = 8'h22;
mem[16'hE065] = 8'hA5;
mem[16'hE066] = 8'h81;
mem[16'hE067] = 8'hD1;
mem[16'hE068] = 8'h9B;
mem[16'hE069] = 8'hD0;
mem[16'hE06A] = 8'h08;
mem[16'hE06B] = 8'hA5;
mem[16'hE06C] = 8'h82;
mem[16'hE06D] = 8'hC8;
mem[16'hE06E] = 8'hD1;
mem[16'hE06F] = 8'h9B;
mem[16'hE070] = 8'hF0;
mem[16'hE071] = 8'h6C;
mem[16'hE072] = 8'h88;
mem[16'hE073] = 8'h18;
mem[16'hE074] = 8'hA5;
mem[16'hE075] = 8'h9B;
mem[16'hE076] = 8'h69;
mem[16'hE077] = 8'h07;
mem[16'hE078] = 8'h90;
mem[16'hE079] = 8'hE1;
mem[16'hE07A] = 8'hE8;
mem[16'hE07B] = 8'hD0;
mem[16'hE07C] = 8'hDC;
mem[16'hE07D] = 8'hC9;
mem[16'hE07E] = 8'h41;
mem[16'hE07F] = 8'h90;
mem[16'hE080] = 8'h05;
mem[16'hE081] = 8'hE9;
mem[16'hE082] = 8'h5B;
mem[16'hE083] = 8'h38;
mem[16'hE084] = 8'hE9;
mem[16'hE085] = 8'hA5;
mem[16'hE086] = 8'h60;
mem[16'hE087] = 8'h68;
mem[16'hE088] = 8'h48;
mem[16'hE089] = 8'hC9;
mem[16'hE08A] = 8'hD7;
mem[16'hE08B] = 8'hD0;
mem[16'hE08C] = 8'h0F;
mem[16'hE08D] = 8'hBA;
mem[16'hE08E] = 8'hBD;
mem[16'hE08F] = 8'h02;
mem[16'hE090] = 8'h01;
mem[16'hE091] = 8'hC9;
mem[16'hE092] = 8'hDE;
mem[16'hE093] = 8'hD0;
mem[16'hE094] = 8'h07;
mem[16'hE095] = 8'hA9;
mem[16'hE096] = 8'h9A;
mem[16'hE097] = 8'hA0;
mem[16'hE098] = 8'hE0;
mem[16'hE099] = 8'h60;
mem[16'hE09A] = 8'h00;
mem[16'hE09B] = 8'h00;
mem[16'hE09C] = 8'hA5;
mem[16'hE09D] = 8'h6B;
mem[16'hE09E] = 8'hA4;
mem[16'hE09F] = 8'h6C;
mem[16'hE0A0] = 8'h85;
mem[16'hE0A1] = 8'h9B;
mem[16'hE0A2] = 8'h84;
mem[16'hE0A3] = 8'h9C;
mem[16'hE0A4] = 8'hA5;
mem[16'hE0A5] = 8'h6D;
mem[16'hE0A6] = 8'hA4;
mem[16'hE0A7] = 8'h6E;
mem[16'hE0A8] = 8'h85;
mem[16'hE0A9] = 8'h96;
mem[16'hE0AA] = 8'h84;
mem[16'hE0AB] = 8'h97;
mem[16'hE0AC] = 8'h18;
mem[16'hE0AD] = 8'h69;
mem[16'hE0AE] = 8'h07;
mem[16'hE0AF] = 8'h90;
mem[16'hE0B0] = 8'h01;
mem[16'hE0B1] = 8'hC8;
mem[16'hE0B2] = 8'h85;
mem[16'hE0B3] = 8'h94;
mem[16'hE0B4] = 8'h84;
mem[16'hE0B5] = 8'h95;
mem[16'hE0B6] = 8'h20;
mem[16'hE0B7] = 8'h93;
mem[16'hE0B8] = 8'hD3;
mem[16'hE0B9] = 8'hA5;
mem[16'hE0BA] = 8'h94;
mem[16'hE0BB] = 8'hA4;
mem[16'hE0BC] = 8'h95;
mem[16'hE0BD] = 8'hC8;
mem[16'hE0BE] = 8'h85;
mem[16'hE0BF] = 8'h6B;
mem[16'hE0C0] = 8'h84;
mem[16'hE0C1] = 8'h6C;
mem[16'hE0C2] = 8'hA0;
mem[16'hE0C3] = 8'h00;
mem[16'hE0C4] = 8'hA5;
mem[16'hE0C5] = 8'h81;
mem[16'hE0C6] = 8'h91;
mem[16'hE0C7] = 8'h9B;
mem[16'hE0C8] = 8'hC8;
mem[16'hE0C9] = 8'hA5;
mem[16'hE0CA] = 8'h82;
mem[16'hE0CB] = 8'h91;
mem[16'hE0CC] = 8'h9B;
mem[16'hE0CD] = 8'hA9;
mem[16'hE0CE] = 8'h00;
mem[16'hE0CF] = 8'hC8;
mem[16'hE0D0] = 8'h91;
mem[16'hE0D1] = 8'h9B;
mem[16'hE0D2] = 8'hC8;
mem[16'hE0D3] = 8'h91;
mem[16'hE0D4] = 8'h9B;
mem[16'hE0D5] = 8'hC8;
mem[16'hE0D6] = 8'h91;
mem[16'hE0D7] = 8'h9B;
mem[16'hE0D8] = 8'hC8;
mem[16'hE0D9] = 8'h91;
mem[16'hE0DA] = 8'h9B;
mem[16'hE0DB] = 8'hC8;
mem[16'hE0DC] = 8'h91;
mem[16'hE0DD] = 8'h9B;
mem[16'hE0DE] = 8'hA5;
mem[16'hE0DF] = 8'h9B;
mem[16'hE0E0] = 8'h18;
mem[16'hE0E1] = 8'h69;
mem[16'hE0E2] = 8'h02;
mem[16'hE0E3] = 8'hA4;
mem[16'hE0E4] = 8'h9C;
mem[16'hE0E5] = 8'h90;
mem[16'hE0E6] = 8'h01;
mem[16'hE0E7] = 8'hC8;
mem[16'hE0E8] = 8'h85;
mem[16'hE0E9] = 8'h83;
mem[16'hE0EA] = 8'h84;
mem[16'hE0EB] = 8'h84;
mem[16'hE0EC] = 8'h60;
mem[16'hE0ED] = 8'hA5;
mem[16'hE0EE] = 8'h0F;
mem[16'hE0EF] = 8'h0A;
mem[16'hE0F0] = 8'h69;
mem[16'hE0F1] = 8'h05;
mem[16'hE0F2] = 8'h65;
mem[16'hE0F3] = 8'h9B;
mem[16'hE0F4] = 8'hA4;
mem[16'hE0F5] = 8'h9C;
mem[16'hE0F6] = 8'h90;
mem[16'hE0F7] = 8'h01;
mem[16'hE0F8] = 8'hC8;
mem[16'hE0F9] = 8'h85;
mem[16'hE0FA] = 8'h94;
mem[16'hE0FB] = 8'h84;
mem[16'hE0FC] = 8'h95;
mem[16'hE0FD] = 8'h60;
mem[16'hE0FE] = 8'h90;
mem[16'hE0FF] = 8'h80;
mem[16'hE100] = 8'h00;
mem[16'hE101] = 8'h00;
mem[16'hE102] = 8'h20;
mem[16'hE103] = 8'hB1;
mem[16'hE104] = 8'h00;
mem[16'hE105] = 8'h20;
mem[16'hE106] = 8'h67;
mem[16'hE107] = 8'hDD;
mem[16'hE108] = 8'hA5;
mem[16'hE109] = 8'hA2;
mem[16'hE10A] = 8'h30;
mem[16'hE10B] = 8'h0D;
mem[16'hE10C] = 8'hA5;
mem[16'hE10D] = 8'h9D;
mem[16'hE10E] = 8'hC9;
mem[16'hE10F] = 8'h90;
mem[16'hE110] = 8'h90;
mem[16'hE111] = 8'h09;
mem[16'hE112] = 8'hA9;
mem[16'hE113] = 8'hFE;
mem[16'hE114] = 8'hA0;
mem[16'hE115] = 8'hE0;
mem[16'hE116] = 8'h20;
mem[16'hE117] = 8'hB2;
mem[16'hE118] = 8'hEB;
mem[16'hE119] = 8'hD0;
mem[16'hE11A] = 8'h7E;
mem[16'hE11B] = 8'h4C;
mem[16'hE11C] = 8'hF2;
mem[16'hE11D] = 8'hEB;
mem[16'hE11E] = 8'hA5;
mem[16'hE11F] = 8'h14;
mem[16'hE120] = 8'hD0;
mem[16'hE121] = 8'h47;
mem[16'hE122] = 8'hA5;
mem[16'hE123] = 8'h10;
mem[16'hE124] = 8'h05;
mem[16'hE125] = 8'h12;
mem[16'hE126] = 8'h48;
mem[16'hE127] = 8'hA5;
mem[16'hE128] = 8'h11;
mem[16'hE129] = 8'h48;
mem[16'hE12A] = 8'hA0;
mem[16'hE12B] = 8'h00;
mem[16'hE12C] = 8'h98;
mem[16'hE12D] = 8'h48;
mem[16'hE12E] = 8'hA5;
mem[16'hE12F] = 8'h82;
mem[16'hE130] = 8'h48;
mem[16'hE131] = 8'hA5;
mem[16'hE132] = 8'h81;
mem[16'hE133] = 8'h48;
mem[16'hE134] = 8'h20;
mem[16'hE135] = 8'h02;
mem[16'hE136] = 8'hE1;
mem[16'hE137] = 8'h68;
mem[16'hE138] = 8'h85;
mem[16'hE139] = 8'h81;
mem[16'hE13A] = 8'h68;
mem[16'hE13B] = 8'h85;
mem[16'hE13C] = 8'h82;
mem[16'hE13D] = 8'h68;
mem[16'hE13E] = 8'hA8;
mem[16'hE13F] = 8'hBA;
mem[16'hE140] = 8'hBD;
mem[16'hE141] = 8'h02;
mem[16'hE142] = 8'h01;
mem[16'hE143] = 8'h48;
mem[16'hE144] = 8'hBD;
mem[16'hE145] = 8'h01;
mem[16'hE146] = 8'h01;
mem[16'hE147] = 8'h48;
mem[16'hE148] = 8'hA5;
mem[16'hE149] = 8'hA0;
mem[16'hE14A] = 8'h9D;
mem[16'hE14B] = 8'h02;
mem[16'hE14C] = 8'h01;
mem[16'hE14D] = 8'hA5;
mem[16'hE14E] = 8'hA1;
mem[16'hE14F] = 8'h9D;
mem[16'hE150] = 8'h01;
mem[16'hE151] = 8'h01;
mem[16'hE152] = 8'hC8;
mem[16'hE153] = 8'h20;
mem[16'hE154] = 8'hB7;
mem[16'hE155] = 8'h00;
mem[16'hE156] = 8'hC9;
mem[16'hE157] = 8'h2C;
mem[16'hE158] = 8'hF0;
mem[16'hE159] = 8'hD2;
mem[16'hE15A] = 8'h84;
mem[16'hE15B] = 8'h0F;
mem[16'hE15C] = 8'h20;
mem[16'hE15D] = 8'hB8;
mem[16'hE15E] = 8'hDE;
mem[16'hE15F] = 8'h68;
mem[16'hE160] = 8'h85;
mem[16'hE161] = 8'h11;
mem[16'hE162] = 8'h68;
mem[16'hE163] = 8'h85;
mem[16'hE164] = 8'h12;
mem[16'hE165] = 8'h29;
mem[16'hE166] = 8'h7F;
mem[16'hE167] = 8'h85;
mem[16'hE168] = 8'h10;
mem[16'hE169] = 8'hA6;
mem[16'hE16A] = 8'h6B;
mem[16'hE16B] = 8'hA5;
mem[16'hE16C] = 8'h6C;
mem[16'hE16D] = 8'h86;
mem[16'hE16E] = 8'h9B;
mem[16'hE16F] = 8'h85;
mem[16'hE170] = 8'h9C;
mem[16'hE171] = 8'hC5;
mem[16'hE172] = 8'h6E;
mem[16'hE173] = 8'hD0;
mem[16'hE174] = 8'h04;
mem[16'hE175] = 8'hE4;
mem[16'hE176] = 8'h6D;
mem[16'hE177] = 8'hF0;
mem[16'hE178] = 8'h3F;
mem[16'hE179] = 8'hA0;
mem[16'hE17A] = 8'h00;
mem[16'hE17B] = 8'hB1;
mem[16'hE17C] = 8'h9B;
mem[16'hE17D] = 8'hC8;
mem[16'hE17E] = 8'hC5;
mem[16'hE17F] = 8'h81;
mem[16'hE180] = 8'hD0;
mem[16'hE181] = 8'h06;
mem[16'hE182] = 8'hA5;
mem[16'hE183] = 8'h82;
mem[16'hE184] = 8'hD1;
mem[16'hE185] = 8'h9B;
mem[16'hE186] = 8'hF0;
mem[16'hE187] = 8'h16;
mem[16'hE188] = 8'hC8;
mem[16'hE189] = 8'hB1;
mem[16'hE18A] = 8'h9B;
mem[16'hE18B] = 8'h18;
mem[16'hE18C] = 8'h65;
mem[16'hE18D] = 8'h9B;
mem[16'hE18E] = 8'hAA;
mem[16'hE18F] = 8'hC8;
mem[16'hE190] = 8'hB1;
mem[16'hE191] = 8'h9B;
mem[16'hE192] = 8'h65;
mem[16'hE193] = 8'h9C;
mem[16'hE194] = 8'h90;
mem[16'hE195] = 8'hD7;
mem[16'hE196] = 8'hA2;
mem[16'hE197] = 8'h6B;
mem[16'hE198] = 8'h2C;
mem[16'hE199] = 8'hA2;
mem[16'hE19A] = 8'h35;
mem[16'hE19B] = 8'h4C;
mem[16'hE19C] = 8'h12;
mem[16'hE19D] = 8'hD4;
mem[16'hE19E] = 8'hA2;
mem[16'hE19F] = 8'h78;
mem[16'hE1A0] = 8'hA5;
mem[16'hE1A1] = 8'h10;
mem[16'hE1A2] = 8'hD0;
mem[16'hE1A3] = 8'hF7;
mem[16'hE1A4] = 8'hA5;
mem[16'hE1A5] = 8'h14;
mem[16'hE1A6] = 8'hF0;
mem[16'hE1A7] = 8'h02;
mem[16'hE1A8] = 8'h38;
mem[16'hE1A9] = 8'h60;
mem[16'hE1AA] = 8'h20;
mem[16'hE1AB] = 8'hED;
mem[16'hE1AC] = 8'hE0;
mem[16'hE1AD] = 8'hA5;
mem[16'hE1AE] = 8'h0F;
mem[16'hE1AF] = 8'hA0;
mem[16'hE1B0] = 8'h04;
mem[16'hE1B1] = 8'hD1;
mem[16'hE1B2] = 8'h9B;
mem[16'hE1B3] = 8'hD0;
mem[16'hE1B4] = 8'hE1;
mem[16'hE1B5] = 8'h4C;
mem[16'hE1B6] = 8'h4B;
mem[16'hE1B7] = 8'hE2;
mem[16'hE1B8] = 8'hA5;
mem[16'hE1B9] = 8'h14;
mem[16'hE1BA] = 8'hF0;
mem[16'hE1BB] = 8'h05;
mem[16'hE1BC] = 8'hA2;
mem[16'hE1BD] = 8'h2A;
mem[16'hE1BE] = 8'h4C;
mem[16'hE1BF] = 8'h12;
mem[16'hE1C0] = 8'hD4;
mem[16'hE1C1] = 8'h20;
mem[16'hE1C2] = 8'hED;
mem[16'hE1C3] = 8'hE0;
mem[16'hE1C4] = 8'h20;
mem[16'hE1C5] = 8'hE3;
mem[16'hE1C6] = 8'hD3;
mem[16'hE1C7] = 8'hA9;
mem[16'hE1C8] = 8'h00;
mem[16'hE1C9] = 8'hA8;
mem[16'hE1CA] = 8'h85;
mem[16'hE1CB] = 8'hAE;
mem[16'hE1CC] = 8'hA2;
mem[16'hE1CD] = 8'h05;
mem[16'hE1CE] = 8'hA5;
mem[16'hE1CF] = 8'h81;
mem[16'hE1D0] = 8'h91;
mem[16'hE1D1] = 8'h9B;
mem[16'hE1D2] = 8'h10;
mem[16'hE1D3] = 8'h01;
mem[16'hE1D4] = 8'hCA;
mem[16'hE1D5] = 8'hC8;
mem[16'hE1D6] = 8'hA5;
mem[16'hE1D7] = 8'h82;
mem[16'hE1D8] = 8'h91;
mem[16'hE1D9] = 8'h9B;
mem[16'hE1DA] = 8'h10;
mem[16'hE1DB] = 8'h02;
mem[16'hE1DC] = 8'hCA;
mem[16'hE1DD] = 8'hCA;
mem[16'hE1DE] = 8'h86;
mem[16'hE1DF] = 8'hAD;
mem[16'hE1E0] = 8'hA5;
mem[16'hE1E1] = 8'h0F;
mem[16'hE1E2] = 8'hC8;
mem[16'hE1E3] = 8'hC8;
mem[16'hE1E4] = 8'hC8;
mem[16'hE1E5] = 8'h91;
mem[16'hE1E6] = 8'h9B;
mem[16'hE1E7] = 8'hA2;
mem[16'hE1E8] = 8'h0B;
mem[16'hE1E9] = 8'hA9;
mem[16'hE1EA] = 8'h00;
mem[16'hE1EB] = 8'h24;
mem[16'hE1EC] = 8'h10;
mem[16'hE1ED] = 8'h50;
mem[16'hE1EE] = 8'h08;
mem[16'hE1EF] = 8'h68;
mem[16'hE1F0] = 8'h18;
mem[16'hE1F1] = 8'h69;
mem[16'hE1F2] = 8'h01;
mem[16'hE1F3] = 8'hAA;
mem[16'hE1F4] = 8'h68;
mem[16'hE1F5] = 8'h69;
mem[16'hE1F6] = 8'h00;
mem[16'hE1F7] = 8'hC8;
mem[16'hE1F8] = 8'h91;
mem[16'hE1F9] = 8'h9B;
mem[16'hE1FA] = 8'hC8;
mem[16'hE1FB] = 8'h8A;
mem[16'hE1FC] = 8'h91;
mem[16'hE1FD] = 8'h9B;
mem[16'hE1FE] = 8'h20;
mem[16'hE1FF] = 8'hAD;
mem[16'hE200] = 8'hE2;
mem[16'hE201] = 8'h86;
mem[16'hE202] = 8'hAD;
mem[16'hE203] = 8'h85;
mem[16'hE204] = 8'hAE;
mem[16'hE205] = 8'hA4;
mem[16'hE206] = 8'h5E;
mem[16'hE207] = 8'hC6;
mem[16'hE208] = 8'h0F;
mem[16'hE209] = 8'hD0;
mem[16'hE20A] = 8'hDC;
mem[16'hE20B] = 8'h65;
mem[16'hE20C] = 8'h95;
mem[16'hE20D] = 8'hB0;
mem[16'hE20E] = 8'h5D;
mem[16'hE20F] = 8'h85;
mem[16'hE210] = 8'h95;
mem[16'hE211] = 8'hA8;
mem[16'hE212] = 8'h8A;
mem[16'hE213] = 8'h65;
mem[16'hE214] = 8'h94;
mem[16'hE215] = 8'h90;
mem[16'hE216] = 8'h03;
mem[16'hE217] = 8'hC8;
mem[16'hE218] = 8'hF0;
mem[16'hE219] = 8'h52;
mem[16'hE21A] = 8'h20;
mem[16'hE21B] = 8'hE3;
mem[16'hE21C] = 8'hD3;
mem[16'hE21D] = 8'h85;
mem[16'hE21E] = 8'h6D;
mem[16'hE21F] = 8'h84;
mem[16'hE220] = 8'h6E;
mem[16'hE221] = 8'hA9;
mem[16'hE222] = 8'h00;
mem[16'hE223] = 8'hE6;
mem[16'hE224] = 8'hAE;
mem[16'hE225] = 8'hA4;
mem[16'hE226] = 8'hAD;
mem[16'hE227] = 8'hF0;
mem[16'hE228] = 8'h05;
mem[16'hE229] = 8'h88;
mem[16'hE22A] = 8'h91;
mem[16'hE22B] = 8'h94;
mem[16'hE22C] = 8'hD0;
mem[16'hE22D] = 8'hFB;
mem[16'hE22E] = 8'hC6;
mem[16'hE22F] = 8'h95;
mem[16'hE230] = 8'hC6;
mem[16'hE231] = 8'hAE;
mem[16'hE232] = 8'hD0;
mem[16'hE233] = 8'hF5;
mem[16'hE234] = 8'hE6;
mem[16'hE235] = 8'h95;
mem[16'hE236] = 8'h38;
mem[16'hE237] = 8'hA5;
mem[16'hE238] = 8'h6D;
mem[16'hE239] = 8'hE5;
mem[16'hE23A] = 8'h9B;
mem[16'hE23B] = 8'hA0;
mem[16'hE23C] = 8'h02;
mem[16'hE23D] = 8'h91;
mem[16'hE23E] = 8'h9B;
mem[16'hE23F] = 8'hA5;
mem[16'hE240] = 8'h6E;
mem[16'hE241] = 8'hC8;
mem[16'hE242] = 8'hE5;
mem[16'hE243] = 8'h9C;
mem[16'hE244] = 8'h91;
mem[16'hE245] = 8'h9B;
mem[16'hE246] = 8'hA5;
mem[16'hE247] = 8'h10;
mem[16'hE248] = 8'hD0;
mem[16'hE249] = 8'h62;
mem[16'hE24A] = 8'hC8;
mem[16'hE24B] = 8'hB1;
mem[16'hE24C] = 8'h9B;
mem[16'hE24D] = 8'h85;
mem[16'hE24E] = 8'h0F;
mem[16'hE24F] = 8'hA9;
mem[16'hE250] = 8'h00;
mem[16'hE251] = 8'h85;
mem[16'hE252] = 8'hAD;
mem[16'hE253] = 8'h85;
mem[16'hE254] = 8'hAE;
mem[16'hE255] = 8'hC8;
mem[16'hE256] = 8'h68;
mem[16'hE257] = 8'hAA;
mem[16'hE258] = 8'h85;
mem[16'hE259] = 8'hA0;
mem[16'hE25A] = 8'h68;
mem[16'hE25B] = 8'h85;
mem[16'hE25C] = 8'hA1;
mem[16'hE25D] = 8'hD1;
mem[16'hE25E] = 8'h9B;
mem[16'hE25F] = 8'h90;
mem[16'hE260] = 8'h0E;
mem[16'hE261] = 8'hD0;
mem[16'hE262] = 8'h06;
mem[16'hE263] = 8'hC8;
mem[16'hE264] = 8'h8A;
mem[16'hE265] = 8'hD1;
mem[16'hE266] = 8'h9B;
mem[16'hE267] = 8'h90;
mem[16'hE268] = 8'h07;
mem[16'hE269] = 8'h4C;
mem[16'hE26A] = 8'h96;
mem[16'hE26B] = 8'hE1;
mem[16'hE26C] = 8'h4C;
mem[16'hE26D] = 8'h10;
mem[16'hE26E] = 8'hD4;
mem[16'hE26F] = 8'hC8;
mem[16'hE270] = 8'hA5;
mem[16'hE271] = 8'hAE;
mem[16'hE272] = 8'h05;
mem[16'hE273] = 8'hAD;
mem[16'hE274] = 8'h18;
mem[16'hE275] = 8'hF0;
mem[16'hE276] = 8'h0A;
mem[16'hE277] = 8'h20;
mem[16'hE278] = 8'hAD;
mem[16'hE279] = 8'hE2;
mem[16'hE27A] = 8'h8A;
mem[16'hE27B] = 8'h65;
mem[16'hE27C] = 8'hA0;
mem[16'hE27D] = 8'hAA;
mem[16'hE27E] = 8'h98;
mem[16'hE27F] = 8'hA4;
mem[16'hE280] = 8'h5E;
mem[16'hE281] = 8'h65;
mem[16'hE282] = 8'hA1;
mem[16'hE283] = 8'h86;
mem[16'hE284] = 8'hAD;
mem[16'hE285] = 8'hC6;
mem[16'hE286] = 8'h0F;
mem[16'hE287] = 8'hD0;
mem[16'hE288] = 8'hCA;
mem[16'hE289] = 8'h85;
mem[16'hE28A] = 8'hAE;
mem[16'hE28B] = 8'hA2;
mem[16'hE28C] = 8'h05;
mem[16'hE28D] = 8'hA5;
mem[16'hE28E] = 8'h81;
mem[16'hE28F] = 8'h10;
mem[16'hE290] = 8'h01;
mem[16'hE291] = 8'hCA;
mem[16'hE292] = 8'hA5;
mem[16'hE293] = 8'h82;
mem[16'hE294] = 8'h10;
mem[16'hE295] = 8'h02;
mem[16'hE296] = 8'hCA;
mem[16'hE297] = 8'hCA;
mem[16'hE298] = 8'h86;
mem[16'hE299] = 8'h64;
mem[16'hE29A] = 8'hA9;
mem[16'hE29B] = 8'h00;
mem[16'hE29C] = 8'h20;
mem[16'hE29D] = 8'hB6;
mem[16'hE29E] = 8'hE2;
mem[16'hE29F] = 8'h8A;
mem[16'hE2A0] = 8'h65;
mem[16'hE2A1] = 8'h94;
mem[16'hE2A2] = 8'h85;
mem[16'hE2A3] = 8'h83;
mem[16'hE2A4] = 8'h98;
mem[16'hE2A5] = 8'h65;
mem[16'hE2A6] = 8'h95;
mem[16'hE2A7] = 8'h85;
mem[16'hE2A8] = 8'h84;
mem[16'hE2A9] = 8'hA8;
mem[16'hE2AA] = 8'hA5;
mem[16'hE2AB] = 8'h83;
mem[16'hE2AC] = 8'h60;
mem[16'hE2AD] = 8'h84;
mem[16'hE2AE] = 8'h5E;
mem[16'hE2AF] = 8'hB1;
mem[16'hE2B0] = 8'h9B;
mem[16'hE2B1] = 8'h85;
mem[16'hE2B2] = 8'h64;
mem[16'hE2B3] = 8'h88;
mem[16'hE2B4] = 8'hB1;
mem[16'hE2B5] = 8'h9B;
mem[16'hE2B6] = 8'h85;
mem[16'hE2B7] = 8'h65;
mem[16'hE2B8] = 8'hA9;
mem[16'hE2B9] = 8'h10;
mem[16'hE2BA] = 8'h85;
mem[16'hE2BB] = 8'h99;
mem[16'hE2BC] = 8'hA2;
mem[16'hE2BD] = 8'h00;
mem[16'hE2BE] = 8'hA0;
mem[16'hE2BF] = 8'h00;
mem[16'hE2C0] = 8'h8A;
mem[16'hE2C1] = 8'h0A;
mem[16'hE2C2] = 8'hAA;
mem[16'hE2C3] = 8'h98;
mem[16'hE2C4] = 8'h2A;
mem[16'hE2C5] = 8'hA8;
mem[16'hE2C6] = 8'hB0;
mem[16'hE2C7] = 8'hA4;
mem[16'hE2C8] = 8'h06;
mem[16'hE2C9] = 8'hAD;
mem[16'hE2CA] = 8'h26;
mem[16'hE2CB] = 8'hAE;
mem[16'hE2CC] = 8'h90;
mem[16'hE2CD] = 8'h0B;
mem[16'hE2CE] = 8'h18;
mem[16'hE2CF] = 8'h8A;
mem[16'hE2D0] = 8'h65;
mem[16'hE2D1] = 8'h64;
mem[16'hE2D2] = 8'hAA;
mem[16'hE2D3] = 8'h98;
mem[16'hE2D4] = 8'h65;
mem[16'hE2D5] = 8'h65;
mem[16'hE2D6] = 8'hA8;
mem[16'hE2D7] = 8'hB0;
mem[16'hE2D8] = 8'h93;
mem[16'hE2D9] = 8'hC6;
mem[16'hE2DA] = 8'h99;
mem[16'hE2DB] = 8'hD0;
mem[16'hE2DC] = 8'hE3;
mem[16'hE2DD] = 8'h60;
mem[16'hE2DE] = 8'hA5;
mem[16'hE2DF] = 8'h11;
mem[16'hE2E0] = 8'hF0;
mem[16'hE2E1] = 8'h03;
mem[16'hE2E2] = 8'h20;
mem[16'hE2E3] = 8'h00;
mem[16'hE2E4] = 8'hE6;
mem[16'hE2E5] = 8'h20;
mem[16'hE2E6] = 8'h84;
mem[16'hE2E7] = 8'hE4;
mem[16'hE2E8] = 8'h38;
mem[16'hE2E9] = 8'hA5;
mem[16'hE2EA] = 8'h6F;
mem[16'hE2EB] = 8'hE5;
mem[16'hE2EC] = 8'h6D;
mem[16'hE2ED] = 8'hA8;
mem[16'hE2EE] = 8'hA5;
mem[16'hE2EF] = 8'h70;
mem[16'hE2F0] = 8'hE5;
mem[16'hE2F1] = 8'h6E;
mem[16'hE2F2] = 8'hA2;
mem[16'hE2F3] = 8'h00;
mem[16'hE2F4] = 8'h86;
mem[16'hE2F5] = 8'h11;
mem[16'hE2F6] = 8'h85;
mem[16'hE2F7] = 8'h9E;
mem[16'hE2F8] = 8'h84;
mem[16'hE2F9] = 8'h9F;
mem[16'hE2FA] = 8'hA2;
mem[16'hE2FB] = 8'h90;
mem[16'hE2FC] = 8'h4C;
mem[16'hE2FD] = 8'h9B;
mem[16'hE2FE] = 8'hEB;
mem[16'hE2FF] = 8'hA4;
mem[16'hE300] = 8'h24;
mem[16'hE301] = 8'hA9;
mem[16'hE302] = 8'h00;
mem[16'hE303] = 8'h38;
mem[16'hE304] = 8'hF0;
mem[16'hE305] = 8'hEC;
mem[16'hE306] = 8'hA6;
mem[16'hE307] = 8'h76;
mem[16'hE308] = 8'hE8;
mem[16'hE309] = 8'hD0;
mem[16'hE30A] = 8'hA1;
mem[16'hE30B] = 8'hA2;
mem[16'hE30C] = 8'h95;
mem[16'hE30D] = 8'h2C;
mem[16'hE30E] = 8'hA2;
mem[16'hE30F] = 8'hE0;
mem[16'hE310] = 8'h4C;
mem[16'hE311] = 8'h12;
mem[16'hE312] = 8'hD4;
mem[16'hE313] = 8'h20;
mem[16'hE314] = 8'h41;
mem[16'hE315] = 8'hE3;
mem[16'hE316] = 8'h20;
mem[16'hE317] = 8'h06;
mem[16'hE318] = 8'hE3;
mem[16'hE319] = 8'h20;
mem[16'hE31A] = 8'hBB;
mem[16'hE31B] = 8'hDE;
mem[16'hE31C] = 8'hA9;
mem[16'hE31D] = 8'h80;
mem[16'hE31E] = 8'h85;
mem[16'hE31F] = 8'h14;
mem[16'hE320] = 8'h20;
mem[16'hE321] = 8'hE3;
mem[16'hE322] = 8'hDF;
mem[16'hE323] = 8'h20;
mem[16'hE324] = 8'h6A;
mem[16'hE325] = 8'hDD;
mem[16'hE326] = 8'h20;
mem[16'hE327] = 8'hB8;
mem[16'hE328] = 8'hDE;
mem[16'hE329] = 8'hA9;
mem[16'hE32A] = 8'hD0;
mem[16'hE32B] = 8'h20;
mem[16'hE32C] = 8'hC0;
mem[16'hE32D] = 8'hDE;
mem[16'hE32E] = 8'h48;
mem[16'hE32F] = 8'hA5;
mem[16'hE330] = 8'h84;
mem[16'hE331] = 8'h48;
mem[16'hE332] = 8'hA5;
mem[16'hE333] = 8'h83;
mem[16'hE334] = 8'h48;
mem[16'hE335] = 8'hA5;
mem[16'hE336] = 8'hB9;
mem[16'hE337] = 8'h48;
mem[16'hE338] = 8'hA5;
mem[16'hE339] = 8'hB8;
mem[16'hE33A] = 8'h48;
mem[16'hE33B] = 8'h20;
mem[16'hE33C] = 8'h95;
mem[16'hE33D] = 8'hD9;
mem[16'hE33E] = 8'h4C;
mem[16'hE33F] = 8'hAF;
mem[16'hE340] = 8'hE3;
mem[16'hE341] = 8'hA9;
mem[16'hE342] = 8'hC2;
mem[16'hE343] = 8'h20;
mem[16'hE344] = 8'hC0;
mem[16'hE345] = 8'hDE;
mem[16'hE346] = 8'h09;
mem[16'hE347] = 8'h80;
mem[16'hE348] = 8'h85;
mem[16'hE349] = 8'h14;
mem[16'hE34A] = 8'h20;
mem[16'hE34B] = 8'hEA;
mem[16'hE34C] = 8'hDF;
mem[16'hE34D] = 8'h85;
mem[16'hE34E] = 8'h8A;
mem[16'hE34F] = 8'h84;
mem[16'hE350] = 8'h8B;
mem[16'hE351] = 8'h4C;
mem[16'hE352] = 8'h6A;
mem[16'hE353] = 8'hDD;
mem[16'hE354] = 8'h20;
mem[16'hE355] = 8'h41;
mem[16'hE356] = 8'hE3;
mem[16'hE357] = 8'hA5;
mem[16'hE358] = 8'h8B;
mem[16'hE359] = 8'h48;
mem[16'hE35A] = 8'hA5;
mem[16'hE35B] = 8'h8A;
mem[16'hE35C] = 8'h48;
mem[16'hE35D] = 8'h20;
mem[16'hE35E] = 8'hB2;
mem[16'hE35F] = 8'hDE;
mem[16'hE360] = 8'h20;
mem[16'hE361] = 8'h6A;
mem[16'hE362] = 8'hDD;
mem[16'hE363] = 8'h68;
mem[16'hE364] = 8'h85;
mem[16'hE365] = 8'h8A;
mem[16'hE366] = 8'h68;
mem[16'hE367] = 8'h85;
mem[16'hE368] = 8'h8B;
mem[16'hE369] = 8'hA0;
mem[16'hE36A] = 8'h02;
mem[16'hE36B] = 8'hB1;
mem[16'hE36C] = 8'h8A;
mem[16'hE36D] = 8'h85;
mem[16'hE36E] = 8'h83;
mem[16'hE36F] = 8'hAA;
mem[16'hE370] = 8'hC8;
mem[16'hE371] = 8'hB1;
mem[16'hE372] = 8'h8A;
mem[16'hE373] = 8'hF0;
mem[16'hE374] = 8'h99;
mem[16'hE375] = 8'h85;
mem[16'hE376] = 8'h84;
mem[16'hE377] = 8'hC8;
mem[16'hE378] = 8'hB1;
mem[16'hE379] = 8'h83;
mem[16'hE37A] = 8'h48;
mem[16'hE37B] = 8'h88;
mem[16'hE37C] = 8'h10;
mem[16'hE37D] = 8'hFA;
mem[16'hE37E] = 8'hA4;
mem[16'hE37F] = 8'h84;
mem[16'hE380] = 8'h20;
mem[16'hE381] = 8'h2B;
mem[16'hE382] = 8'hEB;
mem[16'hE383] = 8'hA5;
mem[16'hE384] = 8'hB9;
mem[16'hE385] = 8'h48;
mem[16'hE386] = 8'hA5;
mem[16'hE387] = 8'hB8;
mem[16'hE388] = 8'h48;
mem[16'hE389] = 8'hB1;
mem[16'hE38A] = 8'h8A;
mem[16'hE38B] = 8'h85;
mem[16'hE38C] = 8'hB8;
mem[16'hE38D] = 8'hC8;
mem[16'hE38E] = 8'hB1;
mem[16'hE38F] = 8'h8A;
mem[16'hE390] = 8'h85;
mem[16'hE391] = 8'hB9;
mem[16'hE392] = 8'hA5;
mem[16'hE393] = 8'h84;
mem[16'hE394] = 8'h48;
mem[16'hE395] = 8'hA5;
mem[16'hE396] = 8'h83;
mem[16'hE397] = 8'h48;
mem[16'hE398] = 8'h20;
mem[16'hE399] = 8'h67;
mem[16'hE39A] = 8'hDD;
mem[16'hE39B] = 8'h68;
mem[16'hE39C] = 8'h85;
mem[16'hE39D] = 8'h8A;
mem[16'hE39E] = 8'h68;
mem[16'hE39F] = 8'h85;
mem[16'hE3A0] = 8'h8B;
mem[16'hE3A1] = 8'h20;
mem[16'hE3A2] = 8'hB7;
mem[16'hE3A3] = 8'h00;
mem[16'hE3A4] = 8'hF0;
mem[16'hE3A5] = 8'h03;
mem[16'hE3A6] = 8'h4C;
mem[16'hE3A7] = 8'hC9;
mem[16'hE3A8] = 8'hDE;
mem[16'hE3A9] = 8'h68;
mem[16'hE3AA] = 8'h85;
mem[16'hE3AB] = 8'hB8;
mem[16'hE3AC] = 8'h68;
mem[16'hE3AD] = 8'h85;
mem[16'hE3AE] = 8'hB9;
mem[16'hE3AF] = 8'hA0;
mem[16'hE3B0] = 8'h00;
mem[16'hE3B1] = 8'h68;
mem[16'hE3B2] = 8'h91;
mem[16'hE3B3] = 8'h8A;
mem[16'hE3B4] = 8'h68;
mem[16'hE3B5] = 8'hC8;
mem[16'hE3B6] = 8'h91;
mem[16'hE3B7] = 8'h8A;
mem[16'hE3B8] = 8'h68;
mem[16'hE3B9] = 8'hC8;
mem[16'hE3BA] = 8'h91;
mem[16'hE3BB] = 8'h8A;
mem[16'hE3BC] = 8'h68;
mem[16'hE3BD] = 8'hC8;
mem[16'hE3BE] = 8'h91;
mem[16'hE3BF] = 8'h8A;
mem[16'hE3C0] = 8'h68;
mem[16'hE3C1] = 8'hC8;
mem[16'hE3C2] = 8'h91;
mem[16'hE3C3] = 8'h8A;
mem[16'hE3C4] = 8'h60;
mem[16'hE3C5] = 8'h20;
mem[16'hE3C6] = 8'h6A;
mem[16'hE3C7] = 8'hDD;
mem[16'hE3C8] = 8'hA0;
mem[16'hE3C9] = 8'h00;
mem[16'hE3CA] = 8'h20;
mem[16'hE3CB] = 8'h36;
mem[16'hE3CC] = 8'hED;
mem[16'hE3CD] = 8'h68;
mem[16'hE3CE] = 8'h68;
mem[16'hE3CF] = 8'hA9;
mem[16'hE3D0] = 8'hFF;
mem[16'hE3D1] = 8'hA0;
mem[16'hE3D2] = 8'h00;
mem[16'hE3D3] = 8'hF0;
mem[16'hE3D4] = 8'h12;
mem[16'hE3D5] = 8'hA6;
mem[16'hE3D6] = 8'hA0;
mem[16'hE3D7] = 8'hA4;
mem[16'hE3D8] = 8'hA1;
mem[16'hE3D9] = 8'h86;
mem[16'hE3DA] = 8'h8C;
mem[16'hE3DB] = 8'h84;
mem[16'hE3DC] = 8'h8D;
mem[16'hE3DD] = 8'h20;
mem[16'hE3DE] = 8'h52;
mem[16'hE3DF] = 8'hE4;
mem[16'hE3E0] = 8'h86;
mem[16'hE3E1] = 8'h9E;
mem[16'hE3E2] = 8'h84;
mem[16'hE3E3] = 8'h9F;
mem[16'hE3E4] = 8'h85;
mem[16'hE3E5] = 8'h9D;
mem[16'hE3E6] = 8'h60;
mem[16'hE3E7] = 8'hA2;
mem[16'hE3E8] = 8'h22;
mem[16'hE3E9] = 8'h86;
mem[16'hE3EA] = 8'h0D;
mem[16'hE3EB] = 8'h86;
mem[16'hE3EC] = 8'h0E;
mem[16'hE3ED] = 8'h85;
mem[16'hE3EE] = 8'hAB;
mem[16'hE3EF] = 8'h84;
mem[16'hE3F0] = 8'hAC;
mem[16'hE3F1] = 8'h85;
mem[16'hE3F2] = 8'h9E;
mem[16'hE3F3] = 8'h84;
mem[16'hE3F4] = 8'h9F;
mem[16'hE3F5] = 8'hA0;
mem[16'hE3F6] = 8'hFF;
mem[16'hE3F7] = 8'hC8;
mem[16'hE3F8] = 8'hB1;
mem[16'hE3F9] = 8'hAB;
mem[16'hE3FA] = 8'hF0;
mem[16'hE3FB] = 8'h0C;
mem[16'hE3FC] = 8'hC5;
mem[16'hE3FD] = 8'h0D;
mem[16'hE3FE] = 8'hF0;
mem[16'hE3FF] = 8'h04;
mem[16'hE400] = 8'hC5;
mem[16'hE401] = 8'h0E;
mem[16'hE402] = 8'hD0;
mem[16'hE403] = 8'hF3;
mem[16'hE404] = 8'hC9;
mem[16'hE405] = 8'h22;
mem[16'hE406] = 8'hF0;
mem[16'hE407] = 8'h01;
mem[16'hE408] = 8'h18;
mem[16'hE409] = 8'h84;
mem[16'hE40A] = 8'h9D;
mem[16'hE40B] = 8'h98;
mem[16'hE40C] = 8'h65;
mem[16'hE40D] = 8'hAB;
mem[16'hE40E] = 8'h85;
mem[16'hE40F] = 8'hAD;
mem[16'hE410] = 8'hA6;
mem[16'hE411] = 8'hAC;
mem[16'hE412] = 8'h90;
mem[16'hE413] = 8'h01;
mem[16'hE414] = 8'hE8;
mem[16'hE415] = 8'h86;
mem[16'hE416] = 8'hAE;
mem[16'hE417] = 8'hA5;
mem[16'hE418] = 8'hAC;
mem[16'hE419] = 8'hF0;
mem[16'hE41A] = 8'h04;
mem[16'hE41B] = 8'hC9;
mem[16'hE41C] = 8'h02;
mem[16'hE41D] = 8'hD0;
mem[16'hE41E] = 8'h0B;
mem[16'hE41F] = 8'h98;
mem[16'hE420] = 8'h20;
mem[16'hE421] = 8'hD5;
mem[16'hE422] = 8'hE3;
mem[16'hE423] = 8'hA6;
mem[16'hE424] = 8'hAB;
mem[16'hE425] = 8'hA4;
mem[16'hE426] = 8'hAC;
mem[16'hE427] = 8'h20;
mem[16'hE428] = 8'hE2;
mem[16'hE429] = 8'hE5;
mem[16'hE42A] = 8'hA6;
mem[16'hE42B] = 8'h52;
mem[16'hE42C] = 8'hE0;
mem[16'hE42D] = 8'h5E;
mem[16'hE42E] = 8'hD0;
mem[16'hE42F] = 8'h05;
mem[16'hE430] = 8'hA2;
mem[16'hE431] = 8'hBF;
mem[16'hE432] = 8'h4C;
mem[16'hE433] = 8'h12;
mem[16'hE434] = 8'hD4;
mem[16'hE435] = 8'hA5;
mem[16'hE436] = 8'h9D;
mem[16'hE437] = 8'h95;
mem[16'hE438] = 8'h00;
mem[16'hE439] = 8'hA5;
mem[16'hE43A] = 8'h9E;
mem[16'hE43B] = 8'h95;
mem[16'hE43C] = 8'h01;
mem[16'hE43D] = 8'hA5;
mem[16'hE43E] = 8'h9F;
mem[16'hE43F] = 8'h95;
mem[16'hE440] = 8'h02;
mem[16'hE441] = 8'hA0;
mem[16'hE442] = 8'h00;
mem[16'hE443] = 8'h86;
mem[16'hE444] = 8'hA0;
mem[16'hE445] = 8'h84;
mem[16'hE446] = 8'hA1;
mem[16'hE447] = 8'h88;
mem[16'hE448] = 8'h84;
mem[16'hE449] = 8'h11;
mem[16'hE44A] = 8'h86;
mem[16'hE44B] = 8'h53;
mem[16'hE44C] = 8'hE8;
mem[16'hE44D] = 8'hE8;
mem[16'hE44E] = 8'hE8;
mem[16'hE44F] = 8'h86;
mem[16'hE450] = 8'h52;
mem[16'hE451] = 8'h60;
mem[16'hE452] = 8'h46;
mem[16'hE453] = 8'h13;
mem[16'hE454] = 8'h48;
mem[16'hE455] = 8'h49;
mem[16'hE456] = 8'hFF;
mem[16'hE457] = 8'h38;
mem[16'hE458] = 8'h65;
mem[16'hE459] = 8'h6F;
mem[16'hE45A] = 8'hA4;
mem[16'hE45B] = 8'h70;
mem[16'hE45C] = 8'hB0;
mem[16'hE45D] = 8'h01;
mem[16'hE45E] = 8'h88;
mem[16'hE45F] = 8'hC4;
mem[16'hE460] = 8'h6E;
mem[16'hE461] = 8'h90;
mem[16'hE462] = 8'h11;
mem[16'hE463] = 8'hD0;
mem[16'hE464] = 8'h04;
mem[16'hE465] = 8'hC5;
mem[16'hE466] = 8'h6D;
mem[16'hE467] = 8'h90;
mem[16'hE468] = 8'h0B;
mem[16'hE469] = 8'h85;
mem[16'hE46A] = 8'h6F;
mem[16'hE46B] = 8'h84;
mem[16'hE46C] = 8'h70;
mem[16'hE46D] = 8'h85;
mem[16'hE46E] = 8'h71;
mem[16'hE46F] = 8'h84;
mem[16'hE470] = 8'h72;
mem[16'hE471] = 8'hAA;
mem[16'hE472] = 8'h68;
mem[16'hE473] = 8'h60;
mem[16'hE474] = 8'hA2;
mem[16'hE475] = 8'h4D;
mem[16'hE476] = 8'hA5;
mem[16'hE477] = 8'h13;
mem[16'hE478] = 8'h30;
mem[16'hE479] = 8'hB8;
mem[16'hE47A] = 8'h20;
mem[16'hE47B] = 8'h84;
mem[16'hE47C] = 8'hE4;
mem[16'hE47D] = 8'hA9;
mem[16'hE47E] = 8'h80;
mem[16'hE47F] = 8'h85;
mem[16'hE480] = 8'h13;
mem[16'hE481] = 8'h68;
mem[16'hE482] = 8'hD0;
mem[16'hE483] = 8'hD0;
mem[16'hE484] = 8'hA6;
mem[16'hE485] = 8'h73;
mem[16'hE486] = 8'hA5;
mem[16'hE487] = 8'h74;
mem[16'hE488] = 8'h86;
mem[16'hE489] = 8'h6F;
mem[16'hE48A] = 8'h85;
mem[16'hE48B] = 8'h70;
mem[16'hE48C] = 8'hA0;
mem[16'hE48D] = 8'h00;
mem[16'hE48E] = 8'h84;
mem[16'hE48F] = 8'h8B;
mem[16'hE490] = 8'hA5;
mem[16'hE491] = 8'h6D;
mem[16'hE492] = 8'hA6;
mem[16'hE493] = 8'h6E;
mem[16'hE494] = 8'h85;
mem[16'hE495] = 8'h9B;
mem[16'hE496] = 8'h86;
mem[16'hE497] = 8'h9C;
mem[16'hE498] = 8'hA9;
mem[16'hE499] = 8'h55;
mem[16'hE49A] = 8'hA2;
mem[16'hE49B] = 8'h00;
mem[16'hE49C] = 8'h85;
mem[16'hE49D] = 8'h5E;
mem[16'hE49E] = 8'h86;
mem[16'hE49F] = 8'h5F;
mem[16'hE4A0] = 8'hC5;
mem[16'hE4A1] = 8'h52;
mem[16'hE4A2] = 8'hF0;
mem[16'hE4A3] = 8'h05;
mem[16'hE4A4] = 8'h20;
mem[16'hE4A5] = 8'h23;
mem[16'hE4A6] = 8'hE5;
mem[16'hE4A7] = 8'hF0;
mem[16'hE4A8] = 8'hF7;
mem[16'hE4A9] = 8'hA9;
mem[16'hE4AA] = 8'h07;
mem[16'hE4AB] = 8'h85;
mem[16'hE4AC] = 8'h8F;
mem[16'hE4AD] = 8'hA5;
mem[16'hE4AE] = 8'h69;
mem[16'hE4AF] = 8'hA6;
mem[16'hE4B0] = 8'h6A;
mem[16'hE4B1] = 8'h85;
mem[16'hE4B2] = 8'h5E;
mem[16'hE4B3] = 8'h86;
mem[16'hE4B4] = 8'h5F;
mem[16'hE4B5] = 8'hE4;
mem[16'hE4B6] = 8'h6C;
mem[16'hE4B7] = 8'hD0;
mem[16'hE4B8] = 8'h04;
mem[16'hE4B9] = 8'hC5;
mem[16'hE4BA] = 8'h6B;
mem[16'hE4BB] = 8'hF0;
mem[16'hE4BC] = 8'h05;
mem[16'hE4BD] = 8'h20;
mem[16'hE4BE] = 8'h19;
mem[16'hE4BF] = 8'hE5;
mem[16'hE4C0] = 8'hF0;
mem[16'hE4C1] = 8'hF3;
mem[16'hE4C2] = 8'h85;
mem[16'hE4C3] = 8'h94;
mem[16'hE4C4] = 8'h86;
mem[16'hE4C5] = 8'h95;
mem[16'hE4C6] = 8'hA9;
mem[16'hE4C7] = 8'h03;
mem[16'hE4C8] = 8'h85;
mem[16'hE4C9] = 8'h8F;
mem[16'hE4CA] = 8'hA5;
mem[16'hE4CB] = 8'h94;
mem[16'hE4CC] = 8'hA6;
mem[16'hE4CD] = 8'h95;
mem[16'hE4CE] = 8'hE4;
mem[16'hE4CF] = 8'h6E;
mem[16'hE4D0] = 8'hD0;
mem[16'hE4D1] = 8'h07;
mem[16'hE4D2] = 8'hC5;
mem[16'hE4D3] = 8'h6D;
mem[16'hE4D4] = 8'hD0;
mem[16'hE4D5] = 8'h03;
mem[16'hE4D6] = 8'h4C;
mem[16'hE4D7] = 8'h62;
mem[16'hE4D8] = 8'hE5;
mem[16'hE4D9] = 8'h85;
mem[16'hE4DA] = 8'h5E;
mem[16'hE4DB] = 8'h86;
mem[16'hE4DC] = 8'h5F;
mem[16'hE4DD] = 8'hA0;
mem[16'hE4DE] = 8'h00;
mem[16'hE4DF] = 8'hB1;
mem[16'hE4E0] = 8'h5E;
mem[16'hE4E1] = 8'hAA;
mem[16'hE4E2] = 8'hC8;
mem[16'hE4E3] = 8'hB1;
mem[16'hE4E4] = 8'h5E;
mem[16'hE4E5] = 8'h08;
mem[16'hE4E6] = 8'hC8;
mem[16'hE4E7] = 8'hB1;
mem[16'hE4E8] = 8'h5E;
mem[16'hE4E9] = 8'h65;
mem[16'hE4EA] = 8'h94;
mem[16'hE4EB] = 8'h85;
mem[16'hE4EC] = 8'h94;
mem[16'hE4ED] = 8'hC8;
mem[16'hE4EE] = 8'hB1;
mem[16'hE4EF] = 8'h5E;
mem[16'hE4F0] = 8'h65;
mem[16'hE4F1] = 8'h95;
mem[16'hE4F2] = 8'h85;
mem[16'hE4F3] = 8'h95;
mem[16'hE4F4] = 8'h28;
mem[16'hE4F5] = 8'h10;
mem[16'hE4F6] = 8'hD3;
mem[16'hE4F7] = 8'h8A;
mem[16'hE4F8] = 8'h30;
mem[16'hE4F9] = 8'hD0;
mem[16'hE4FA] = 8'hC8;
mem[16'hE4FB] = 8'hB1;
mem[16'hE4FC] = 8'h5E;
mem[16'hE4FD] = 8'hA0;
mem[16'hE4FE] = 8'h00;
mem[16'hE4FF] = 8'h0A;
mem[16'hE500] = 8'h69;
mem[16'hE501] = 8'h05;
mem[16'hE502] = 8'h65;
mem[16'hE503] = 8'h5E;
mem[16'hE504] = 8'h85;
mem[16'hE505] = 8'h5E;
mem[16'hE506] = 8'h90;
mem[16'hE507] = 8'h02;
mem[16'hE508] = 8'hE6;
mem[16'hE509] = 8'h5F;
mem[16'hE50A] = 8'hA6;
mem[16'hE50B] = 8'h5F;
mem[16'hE50C] = 8'hE4;
mem[16'hE50D] = 8'h95;
mem[16'hE50E] = 8'hD0;
mem[16'hE50F] = 8'h04;
mem[16'hE510] = 8'hC5;
mem[16'hE511] = 8'h94;
mem[16'hE512] = 8'hF0;
mem[16'hE513] = 8'hBA;
mem[16'hE514] = 8'h20;
mem[16'hE515] = 8'h23;
mem[16'hE516] = 8'hE5;
mem[16'hE517] = 8'hF0;
mem[16'hE518] = 8'hF3;
mem[16'hE519] = 8'hB1;
mem[16'hE51A] = 8'h5E;
mem[16'hE51B] = 8'h30;
mem[16'hE51C] = 8'h35;
mem[16'hE51D] = 8'hC8;
mem[16'hE51E] = 8'hB1;
mem[16'hE51F] = 8'h5E;
mem[16'hE520] = 8'h10;
mem[16'hE521] = 8'h30;
mem[16'hE522] = 8'hC8;
mem[16'hE523] = 8'hB1;
mem[16'hE524] = 8'h5E;
mem[16'hE525] = 8'hF0;
mem[16'hE526] = 8'h2B;
mem[16'hE527] = 8'hC8;
mem[16'hE528] = 8'hB1;
mem[16'hE529] = 8'h5E;
mem[16'hE52A] = 8'hAA;
mem[16'hE52B] = 8'hC8;
mem[16'hE52C] = 8'hB1;
mem[16'hE52D] = 8'h5E;
mem[16'hE52E] = 8'hC5;
mem[16'hE52F] = 8'h70;
mem[16'hE530] = 8'h90;
mem[16'hE531] = 8'h06;
mem[16'hE532] = 8'hD0;
mem[16'hE533] = 8'h1E;
mem[16'hE534] = 8'hE4;
mem[16'hE535] = 8'h6F;
mem[16'hE536] = 8'hB0;
mem[16'hE537] = 8'h1A;
mem[16'hE538] = 8'hC5;
mem[16'hE539] = 8'h9C;
mem[16'hE53A] = 8'h90;
mem[16'hE53B] = 8'h16;
mem[16'hE53C] = 8'hD0;
mem[16'hE53D] = 8'h04;
mem[16'hE53E] = 8'hE4;
mem[16'hE53F] = 8'h9B;
mem[16'hE540] = 8'h90;
mem[16'hE541] = 8'h10;
mem[16'hE542] = 8'h86;
mem[16'hE543] = 8'h9B;
mem[16'hE544] = 8'h85;
mem[16'hE545] = 8'h9C;
mem[16'hE546] = 8'hA5;
mem[16'hE547] = 8'h5E;
mem[16'hE548] = 8'hA6;
mem[16'hE549] = 8'h5F;
mem[16'hE54A] = 8'h85;
mem[16'hE54B] = 8'h8A;
mem[16'hE54C] = 8'h86;
mem[16'hE54D] = 8'h8B;
mem[16'hE54E] = 8'hA5;
mem[16'hE54F] = 8'h8F;
mem[16'hE550] = 8'h85;
mem[16'hE551] = 8'h91;
mem[16'hE552] = 8'hA5;
mem[16'hE553] = 8'h8F;
mem[16'hE554] = 8'h18;
mem[16'hE555] = 8'h65;
mem[16'hE556] = 8'h5E;
mem[16'hE557] = 8'h85;
mem[16'hE558] = 8'h5E;
mem[16'hE559] = 8'h90;
mem[16'hE55A] = 8'h02;
mem[16'hE55B] = 8'hE6;
mem[16'hE55C] = 8'h5F;
mem[16'hE55D] = 8'hA6;
mem[16'hE55E] = 8'h5F;
mem[16'hE55F] = 8'hA0;
mem[16'hE560] = 8'h00;
mem[16'hE561] = 8'h60;
mem[16'hE562] = 8'hA6;
mem[16'hE563] = 8'h8B;
mem[16'hE564] = 8'hF0;
mem[16'hE565] = 8'hF7;
mem[16'hE566] = 8'hA5;
mem[16'hE567] = 8'h91;
mem[16'hE568] = 8'h29;
mem[16'hE569] = 8'h04;
mem[16'hE56A] = 8'h4A;
mem[16'hE56B] = 8'hA8;
mem[16'hE56C] = 8'h85;
mem[16'hE56D] = 8'h91;
mem[16'hE56E] = 8'hB1;
mem[16'hE56F] = 8'h8A;
mem[16'hE570] = 8'h65;
mem[16'hE571] = 8'h9B;
mem[16'hE572] = 8'h85;
mem[16'hE573] = 8'h96;
mem[16'hE574] = 8'hA5;
mem[16'hE575] = 8'h9C;
mem[16'hE576] = 8'h69;
mem[16'hE577] = 8'h00;
mem[16'hE578] = 8'h85;
mem[16'hE579] = 8'h97;
mem[16'hE57A] = 8'hA5;
mem[16'hE57B] = 8'h6F;
mem[16'hE57C] = 8'hA6;
mem[16'hE57D] = 8'h70;
mem[16'hE57E] = 8'h85;
mem[16'hE57F] = 8'h94;
mem[16'hE580] = 8'h86;
mem[16'hE581] = 8'h95;
mem[16'hE582] = 8'h20;
mem[16'hE583] = 8'h9A;
mem[16'hE584] = 8'hD3;
mem[16'hE585] = 8'hA4;
mem[16'hE586] = 8'h91;
mem[16'hE587] = 8'hC8;
mem[16'hE588] = 8'hA5;
mem[16'hE589] = 8'h94;
mem[16'hE58A] = 8'h91;
mem[16'hE58B] = 8'h8A;
mem[16'hE58C] = 8'hAA;
mem[16'hE58D] = 8'hE6;
mem[16'hE58E] = 8'h95;
mem[16'hE58F] = 8'hA5;
mem[16'hE590] = 8'h95;
mem[16'hE591] = 8'hC8;
mem[16'hE592] = 8'h91;
mem[16'hE593] = 8'h8A;
mem[16'hE594] = 8'h4C;
mem[16'hE595] = 8'h88;
mem[16'hE596] = 8'hE4;
mem[16'hE597] = 8'hA5;
mem[16'hE598] = 8'hA1;
mem[16'hE599] = 8'h48;
mem[16'hE59A] = 8'hA5;
mem[16'hE59B] = 8'hA0;
mem[16'hE59C] = 8'h48;
mem[16'hE59D] = 8'h20;
mem[16'hE59E] = 8'h60;
mem[16'hE59F] = 8'hDE;
mem[16'hE5A0] = 8'h20;
mem[16'hE5A1] = 8'h6C;
mem[16'hE5A2] = 8'hDD;
mem[16'hE5A3] = 8'h68;
mem[16'hE5A4] = 8'h85;
mem[16'hE5A5] = 8'hAB;
mem[16'hE5A6] = 8'h68;
mem[16'hE5A7] = 8'h85;
mem[16'hE5A8] = 8'hAC;
mem[16'hE5A9] = 8'hA0;
mem[16'hE5AA] = 8'h00;
mem[16'hE5AB] = 8'hB1;
mem[16'hE5AC] = 8'hAB;
mem[16'hE5AD] = 8'h18;
mem[16'hE5AE] = 8'h71;
mem[16'hE5AF] = 8'hA0;
mem[16'hE5B0] = 8'h90;
mem[16'hE5B1] = 8'h05;
mem[16'hE5B2] = 8'hA2;
mem[16'hE5B3] = 8'hB0;
mem[16'hE5B4] = 8'h4C;
mem[16'hE5B5] = 8'h12;
mem[16'hE5B6] = 8'hD4;
mem[16'hE5B7] = 8'h20;
mem[16'hE5B8] = 8'hD5;
mem[16'hE5B9] = 8'hE3;
mem[16'hE5BA] = 8'h20;
mem[16'hE5BB] = 8'hD4;
mem[16'hE5BC] = 8'hE5;
mem[16'hE5BD] = 8'hA5;
mem[16'hE5BE] = 8'h8C;
mem[16'hE5BF] = 8'hA4;
mem[16'hE5C0] = 8'h8D;
mem[16'hE5C1] = 8'h20;
mem[16'hE5C2] = 8'h04;
mem[16'hE5C3] = 8'hE6;
mem[16'hE5C4] = 8'h20;
mem[16'hE5C5] = 8'hE6;
mem[16'hE5C6] = 8'hE5;
mem[16'hE5C7] = 8'hA5;
mem[16'hE5C8] = 8'hAB;
mem[16'hE5C9] = 8'hA4;
mem[16'hE5CA] = 8'hAC;
mem[16'hE5CB] = 8'h20;
mem[16'hE5CC] = 8'h04;
mem[16'hE5CD] = 8'hE6;
mem[16'hE5CE] = 8'h20;
mem[16'hE5CF] = 8'h2A;
mem[16'hE5D0] = 8'hE4;
mem[16'hE5D1] = 8'h4C;
mem[16'hE5D2] = 8'h95;
mem[16'hE5D3] = 8'hDD;
mem[16'hE5D4] = 8'hA0;
mem[16'hE5D5] = 8'h00;
mem[16'hE5D6] = 8'hB1;
mem[16'hE5D7] = 8'hAB;
mem[16'hE5D8] = 8'h48;
mem[16'hE5D9] = 8'hC8;
mem[16'hE5DA] = 8'hB1;
mem[16'hE5DB] = 8'hAB;
mem[16'hE5DC] = 8'hAA;
mem[16'hE5DD] = 8'hC8;
mem[16'hE5DE] = 8'hB1;
mem[16'hE5DF] = 8'hAB;
mem[16'hE5E0] = 8'hA8;
mem[16'hE5E1] = 8'h68;
mem[16'hE5E2] = 8'h86;
mem[16'hE5E3] = 8'h5E;
mem[16'hE5E4] = 8'h84;
mem[16'hE5E5] = 8'h5F;
mem[16'hE5E6] = 8'hA8;
mem[16'hE5E7] = 8'hF0;
mem[16'hE5E8] = 8'h0A;
mem[16'hE5E9] = 8'h48;
mem[16'hE5EA] = 8'h88;
mem[16'hE5EB] = 8'hB1;
mem[16'hE5EC] = 8'h5E;
mem[16'hE5ED] = 8'h91;
mem[16'hE5EE] = 8'h71;
mem[16'hE5EF] = 8'h98;
mem[16'hE5F0] = 8'hD0;
mem[16'hE5F1] = 8'hF8;
mem[16'hE5F2] = 8'h68;
mem[16'hE5F3] = 8'h18;
mem[16'hE5F4] = 8'h65;
mem[16'hE5F5] = 8'h71;
mem[16'hE5F6] = 8'h85;
mem[16'hE5F7] = 8'h71;
mem[16'hE5F8] = 8'h90;
mem[16'hE5F9] = 8'h02;
mem[16'hE5FA] = 8'hE6;
mem[16'hE5FB] = 8'h72;
mem[16'hE5FC] = 8'h60;
mem[16'hE5FD] = 8'h20;
mem[16'hE5FE] = 8'h6C;
mem[16'hE5FF] = 8'hDD;
mem[16'hE600] = 8'hA5;
mem[16'hE601] = 8'hA0;
mem[16'hE602] = 8'hA4;
mem[16'hE603] = 8'hA1;
mem[16'hE604] = 8'h85;
mem[16'hE605] = 8'h5E;
mem[16'hE606] = 8'h84;
mem[16'hE607] = 8'h5F;
mem[16'hE608] = 8'h20;
mem[16'hE609] = 8'h35;
mem[16'hE60A] = 8'hE6;
mem[16'hE60B] = 8'h08;
mem[16'hE60C] = 8'hA0;
mem[16'hE60D] = 8'h00;
mem[16'hE60E] = 8'hB1;
mem[16'hE60F] = 8'h5E;
mem[16'hE610] = 8'h48;
mem[16'hE611] = 8'hC8;
mem[16'hE612] = 8'hB1;
mem[16'hE613] = 8'h5E;
mem[16'hE614] = 8'hAA;
mem[16'hE615] = 8'hC8;
mem[16'hE616] = 8'hB1;
mem[16'hE617] = 8'h5E;
mem[16'hE618] = 8'hA8;
mem[16'hE619] = 8'h68;
mem[16'hE61A] = 8'h28;
mem[16'hE61B] = 8'hD0;
mem[16'hE61C] = 8'h13;
mem[16'hE61D] = 8'hC4;
mem[16'hE61E] = 8'h70;
mem[16'hE61F] = 8'hD0;
mem[16'hE620] = 8'h0F;
mem[16'hE621] = 8'hE4;
mem[16'hE622] = 8'h6F;
mem[16'hE623] = 8'hD0;
mem[16'hE624] = 8'h0B;
mem[16'hE625] = 8'h48;
mem[16'hE626] = 8'h18;
mem[16'hE627] = 8'h65;
mem[16'hE628] = 8'h6F;
mem[16'hE629] = 8'h85;
mem[16'hE62A] = 8'h6F;
mem[16'hE62B] = 8'h90;
mem[16'hE62C] = 8'h02;
mem[16'hE62D] = 8'hE6;
mem[16'hE62E] = 8'h70;
mem[16'hE62F] = 8'h68;
mem[16'hE630] = 8'h86;
mem[16'hE631] = 8'h5E;
mem[16'hE632] = 8'h84;
mem[16'hE633] = 8'h5F;
mem[16'hE634] = 8'h60;
mem[16'hE635] = 8'hC4;
mem[16'hE636] = 8'h54;
mem[16'hE637] = 8'hD0;
mem[16'hE638] = 8'h0C;
mem[16'hE639] = 8'hC5;
mem[16'hE63A] = 8'h53;
mem[16'hE63B] = 8'hD0;
mem[16'hE63C] = 8'h08;
mem[16'hE63D] = 8'h85;
mem[16'hE63E] = 8'h52;
mem[16'hE63F] = 8'hE9;
mem[16'hE640] = 8'h03;
mem[16'hE641] = 8'h85;
mem[16'hE642] = 8'h53;
mem[16'hE643] = 8'hA0;
mem[16'hE644] = 8'h00;
mem[16'hE645] = 8'h60;
mem[16'hE646] = 8'h20;
mem[16'hE647] = 8'hFB;
mem[16'hE648] = 8'hE6;
mem[16'hE649] = 8'h8A;
mem[16'hE64A] = 8'h48;
mem[16'hE64B] = 8'hA9;
mem[16'hE64C] = 8'h01;
mem[16'hE64D] = 8'h20;
mem[16'hE64E] = 8'hDD;
mem[16'hE64F] = 8'hE3;
mem[16'hE650] = 8'h68;
mem[16'hE651] = 8'hA0;
mem[16'hE652] = 8'h00;
mem[16'hE653] = 8'h91;
mem[16'hE654] = 8'h9E;
mem[16'hE655] = 8'h68;
mem[16'hE656] = 8'h68;
mem[16'hE657] = 8'h4C;
mem[16'hE658] = 8'h2A;
mem[16'hE659] = 8'hE4;
mem[16'hE65A] = 8'h20;
mem[16'hE65B] = 8'hB9;
mem[16'hE65C] = 8'hE6;
mem[16'hE65D] = 8'hD1;
mem[16'hE65E] = 8'h8C;
mem[16'hE65F] = 8'h98;
mem[16'hE660] = 8'h90;
mem[16'hE661] = 8'h04;
mem[16'hE662] = 8'hB1;
mem[16'hE663] = 8'h8C;
mem[16'hE664] = 8'hAA;
mem[16'hE665] = 8'h98;
mem[16'hE666] = 8'h48;
mem[16'hE667] = 8'h8A;
mem[16'hE668] = 8'h48;
mem[16'hE669] = 8'h20;
mem[16'hE66A] = 8'hDD;
mem[16'hE66B] = 8'hE3;
mem[16'hE66C] = 8'hA5;
mem[16'hE66D] = 8'h8C;
mem[16'hE66E] = 8'hA4;
mem[16'hE66F] = 8'h8D;
mem[16'hE670] = 8'h20;
mem[16'hE671] = 8'h04;
mem[16'hE672] = 8'hE6;
mem[16'hE673] = 8'h68;
mem[16'hE674] = 8'hA8;
mem[16'hE675] = 8'h68;
mem[16'hE676] = 8'h18;
mem[16'hE677] = 8'h65;
mem[16'hE678] = 8'h5E;
mem[16'hE679] = 8'h85;
mem[16'hE67A] = 8'h5E;
mem[16'hE67B] = 8'h90;
mem[16'hE67C] = 8'h02;
mem[16'hE67D] = 8'hE6;
mem[16'hE67E] = 8'h5F;
mem[16'hE67F] = 8'h98;
mem[16'hE680] = 8'h20;
mem[16'hE681] = 8'hE6;
mem[16'hE682] = 8'hE5;
mem[16'hE683] = 8'h4C;
mem[16'hE684] = 8'h2A;
mem[16'hE685] = 8'hE4;
mem[16'hE686] = 8'h20;
mem[16'hE687] = 8'hB9;
mem[16'hE688] = 8'hE6;
mem[16'hE689] = 8'h18;
mem[16'hE68A] = 8'hF1;
mem[16'hE68B] = 8'h8C;
mem[16'hE68C] = 8'h49;
mem[16'hE68D] = 8'hFF;
mem[16'hE68E] = 8'h4C;
mem[16'hE68F] = 8'h60;
mem[16'hE690] = 8'hE6;
mem[16'hE691] = 8'hA9;
mem[16'hE692] = 8'hFF;
mem[16'hE693] = 8'h85;
mem[16'hE694] = 8'hA1;
mem[16'hE695] = 8'h20;
mem[16'hE696] = 8'hB7;
mem[16'hE697] = 8'h00;
mem[16'hE698] = 8'hC9;
mem[16'hE699] = 8'h29;
mem[16'hE69A] = 8'hF0;
mem[16'hE69B] = 8'h06;
mem[16'hE69C] = 8'h20;
mem[16'hE69D] = 8'hBE;
mem[16'hE69E] = 8'hDE;
mem[16'hE69F] = 8'h20;
mem[16'hE6A0] = 8'hF8;
mem[16'hE6A1] = 8'hE6;
mem[16'hE6A2] = 8'h20;
mem[16'hE6A3] = 8'hB9;
mem[16'hE6A4] = 8'hE6;
mem[16'hE6A5] = 8'hCA;
mem[16'hE6A6] = 8'h8A;
mem[16'hE6A7] = 8'h48;
mem[16'hE6A8] = 8'h18;
mem[16'hE6A9] = 8'hA2;
mem[16'hE6AA] = 8'h00;
mem[16'hE6AB] = 8'hF1;
mem[16'hE6AC] = 8'h8C;
mem[16'hE6AD] = 8'hB0;
mem[16'hE6AE] = 8'hB8;
mem[16'hE6AF] = 8'h49;
mem[16'hE6B0] = 8'hFF;
mem[16'hE6B1] = 8'hC5;
mem[16'hE6B2] = 8'hA1;
mem[16'hE6B3] = 8'h90;
mem[16'hE6B4] = 8'hB3;
mem[16'hE6B5] = 8'hA5;
mem[16'hE6B6] = 8'hA1;
mem[16'hE6B7] = 8'hB0;
mem[16'hE6B8] = 8'hAF;
mem[16'hE6B9] = 8'h20;
mem[16'hE6BA] = 8'hB8;
mem[16'hE6BB] = 8'hDE;
mem[16'hE6BC] = 8'h68;
mem[16'hE6BD] = 8'hA8;
mem[16'hE6BE] = 8'h68;
mem[16'hE6BF] = 8'h85;
mem[16'hE6C0] = 8'h91;
mem[16'hE6C1] = 8'h68;
mem[16'hE6C2] = 8'h68;
mem[16'hE6C3] = 8'h68;
mem[16'hE6C4] = 8'hAA;
mem[16'hE6C5] = 8'h68;
mem[16'hE6C6] = 8'h85;
mem[16'hE6C7] = 8'h8C;
mem[16'hE6C8] = 8'h68;
mem[16'hE6C9] = 8'h85;
mem[16'hE6CA] = 8'h8D;
mem[16'hE6CB] = 8'hA5;
mem[16'hE6CC] = 8'h91;
mem[16'hE6CD] = 8'h48;
mem[16'hE6CE] = 8'h98;
mem[16'hE6CF] = 8'h48;
mem[16'hE6D0] = 8'hA0;
mem[16'hE6D1] = 8'h00;
mem[16'hE6D2] = 8'h8A;
mem[16'hE6D3] = 8'hF0;
mem[16'hE6D4] = 8'h1D;
mem[16'hE6D5] = 8'h60;
mem[16'hE6D6] = 8'h20;
mem[16'hE6D7] = 8'hDC;
mem[16'hE6D8] = 8'hE6;
mem[16'hE6D9] = 8'h4C;
mem[16'hE6DA] = 8'h01;
mem[16'hE6DB] = 8'hE3;
mem[16'hE6DC] = 8'h20;
mem[16'hE6DD] = 8'hFD;
mem[16'hE6DE] = 8'hE5;
mem[16'hE6DF] = 8'hA2;
mem[16'hE6E0] = 8'h00;
mem[16'hE6E1] = 8'h86;
mem[16'hE6E2] = 8'h11;
mem[16'hE6E3] = 8'hA8;
mem[16'hE6E4] = 8'h60;
mem[16'hE6E5] = 8'h20;
mem[16'hE6E6] = 8'hDC;
mem[16'hE6E7] = 8'hE6;
mem[16'hE6E8] = 8'hF0;
mem[16'hE6E9] = 8'h08;
mem[16'hE6EA] = 8'hA0;
mem[16'hE6EB] = 8'h00;
mem[16'hE6EC] = 8'hB1;
mem[16'hE6ED] = 8'h5E;
mem[16'hE6EE] = 8'hA8;
mem[16'hE6EF] = 8'h4C;
mem[16'hE6F0] = 8'h01;
mem[16'hE6F1] = 8'hE3;
mem[16'hE6F2] = 8'h4C;
mem[16'hE6F3] = 8'h99;
mem[16'hE6F4] = 8'hE1;
mem[16'hE6F5] = 8'h20;
mem[16'hE6F6] = 8'hB1;
mem[16'hE6F7] = 8'h00;
mem[16'hE6F8] = 8'h20;
mem[16'hE6F9] = 8'h67;
mem[16'hE6FA] = 8'hDD;
mem[16'hE6FB] = 8'h20;
mem[16'hE6FC] = 8'h08;
mem[16'hE6FD] = 8'hE1;
mem[16'hE6FE] = 8'hA6;
mem[16'hE6FF] = 8'hA0;
mem[16'hE700] = 8'hD0;
mem[16'hE701] = 8'hF0;
mem[16'hE702] = 8'hA6;
mem[16'hE703] = 8'hA1;
mem[16'hE704] = 8'h4C;
mem[16'hE705] = 8'hB7;
mem[16'hE706] = 8'h00;
mem[16'hE707] = 8'h20;
mem[16'hE708] = 8'hDC;
mem[16'hE709] = 8'hE6;
mem[16'hE70A] = 8'hD0;
mem[16'hE70B] = 8'h03;
mem[16'hE70C] = 8'h4C;
mem[16'hE70D] = 8'h4E;
mem[16'hE70E] = 8'hE8;
mem[16'hE70F] = 8'hA6;
mem[16'hE710] = 8'hB8;
mem[16'hE711] = 8'hA4;
mem[16'hE712] = 8'hB9;
mem[16'hE713] = 8'h86;
mem[16'hE714] = 8'hAD;
mem[16'hE715] = 8'h84;
mem[16'hE716] = 8'hAE;
mem[16'hE717] = 8'hA6;
mem[16'hE718] = 8'h5E;
mem[16'hE719] = 8'h86;
mem[16'hE71A] = 8'hB8;
mem[16'hE71B] = 8'h18;
mem[16'hE71C] = 8'h65;
mem[16'hE71D] = 8'h5E;
mem[16'hE71E] = 8'h85;
mem[16'hE71F] = 8'h60;
mem[16'hE720] = 8'hA6;
mem[16'hE721] = 8'h5F;
mem[16'hE722] = 8'h86;
mem[16'hE723] = 8'hB9;
mem[16'hE724] = 8'h90;
mem[16'hE725] = 8'h01;
mem[16'hE726] = 8'hE8;
mem[16'hE727] = 8'h86;
mem[16'hE728] = 8'h61;
mem[16'hE729] = 8'hA0;
mem[16'hE72A] = 8'h00;
mem[16'hE72B] = 8'hB1;
mem[16'hE72C] = 8'h60;
mem[16'hE72D] = 8'h48;
mem[16'hE72E] = 8'hA9;
mem[16'hE72F] = 8'h00;
mem[16'hE730] = 8'h91;
mem[16'hE731] = 8'h60;
mem[16'hE732] = 8'h20;
mem[16'hE733] = 8'hB7;
mem[16'hE734] = 8'h00;
mem[16'hE735] = 8'h20;
mem[16'hE736] = 8'h4A;
mem[16'hE737] = 8'hEC;
mem[16'hE738] = 8'h68;
mem[16'hE739] = 8'hA0;
mem[16'hE73A] = 8'h00;
mem[16'hE73B] = 8'h91;
mem[16'hE73C] = 8'h60;
mem[16'hE73D] = 8'hA6;
mem[16'hE73E] = 8'hAD;
mem[16'hE73F] = 8'hA4;
mem[16'hE740] = 8'hAE;
mem[16'hE741] = 8'h86;
mem[16'hE742] = 8'hB8;
mem[16'hE743] = 8'h84;
mem[16'hE744] = 8'hB9;
mem[16'hE745] = 8'h60;
mem[16'hE746] = 8'h20;
mem[16'hE747] = 8'h67;
mem[16'hE748] = 8'hDD;
mem[16'hE749] = 8'h20;
mem[16'hE74A] = 8'h52;
mem[16'hE74B] = 8'hE7;
mem[16'hE74C] = 8'h20;
mem[16'hE74D] = 8'hBE;
mem[16'hE74E] = 8'hDE;
mem[16'hE74F] = 8'h4C;
mem[16'hE750] = 8'hF8;
mem[16'hE751] = 8'hE6;
mem[16'hE752] = 8'hA5;
mem[16'hE753] = 8'h9D;
mem[16'hE754] = 8'hC9;
mem[16'hE755] = 8'h91;
mem[16'hE756] = 8'hB0;
mem[16'hE757] = 8'h9A;
mem[16'hE758] = 8'h20;
mem[16'hE759] = 8'hF2;
mem[16'hE75A] = 8'hEB;
mem[16'hE75B] = 8'hA5;
mem[16'hE75C] = 8'hA0;
mem[16'hE75D] = 8'hA4;
mem[16'hE75E] = 8'hA1;
mem[16'hE75F] = 8'h84;
mem[16'hE760] = 8'h50;
mem[16'hE761] = 8'h85;
mem[16'hE762] = 8'h51;
mem[16'hE763] = 8'h60;
mem[16'hE764] = 8'hA5;
mem[16'hE765] = 8'h50;
mem[16'hE766] = 8'h48;
mem[16'hE767] = 8'hA5;
mem[16'hE768] = 8'h51;
mem[16'hE769] = 8'h48;
mem[16'hE76A] = 8'h20;
mem[16'hE76B] = 8'h52;
mem[16'hE76C] = 8'hE7;
mem[16'hE76D] = 8'hA0;
mem[16'hE76E] = 8'h00;
mem[16'hE76F] = 8'hB1;
mem[16'hE770] = 8'h50;
mem[16'hE771] = 8'hA8;
mem[16'hE772] = 8'h68;
mem[16'hE773] = 8'h85;
mem[16'hE774] = 8'h51;
mem[16'hE775] = 8'h68;
mem[16'hE776] = 8'h85;
mem[16'hE777] = 8'h50;
mem[16'hE778] = 8'h4C;
mem[16'hE779] = 8'h01;
mem[16'hE77A] = 8'hE3;
mem[16'hE77B] = 8'h20;
mem[16'hE77C] = 8'h46;
mem[16'hE77D] = 8'hE7;
mem[16'hE77E] = 8'h8A;
mem[16'hE77F] = 8'hA0;
mem[16'hE780] = 8'h00;
mem[16'hE781] = 8'h91;
mem[16'hE782] = 8'h50;
mem[16'hE783] = 8'h60;
mem[16'hE784] = 8'h20;
mem[16'hE785] = 8'h46;
mem[16'hE786] = 8'hE7;
mem[16'hE787] = 8'h86;
mem[16'hE788] = 8'h85;
mem[16'hE789] = 8'hA2;
mem[16'hE78A] = 8'h00;
mem[16'hE78B] = 8'h20;
mem[16'hE78C] = 8'hB7;
mem[16'hE78D] = 8'h00;
mem[16'hE78E] = 8'hF0;
mem[16'hE78F] = 8'h03;
mem[16'hE790] = 8'h20;
mem[16'hE791] = 8'h4C;
mem[16'hE792] = 8'hE7;
mem[16'hE793] = 8'h86;
mem[16'hE794] = 8'h86;
mem[16'hE795] = 8'hA0;
mem[16'hE796] = 8'h00;
mem[16'hE797] = 8'hB1;
mem[16'hE798] = 8'h50;
mem[16'hE799] = 8'h45;
mem[16'hE79A] = 8'h86;
mem[16'hE79B] = 8'h25;
mem[16'hE79C] = 8'h85;
mem[16'hE79D] = 8'hF0;
mem[16'hE79E] = 8'hF8;
mem[16'hE79F] = 8'h60;
mem[16'hE7A0] = 8'hA9;
mem[16'hE7A1] = 8'h64;
mem[16'hE7A2] = 8'hA0;
mem[16'hE7A3] = 8'hEE;
mem[16'hE7A4] = 8'h4C;
mem[16'hE7A5] = 8'hBE;
mem[16'hE7A6] = 8'hE7;
mem[16'hE7A7] = 8'h20;
mem[16'hE7A8] = 8'hE3;
mem[16'hE7A9] = 8'hE9;
mem[16'hE7AA] = 8'hA5;
mem[16'hE7AB] = 8'hA2;
mem[16'hE7AC] = 8'h49;
mem[16'hE7AD] = 8'hFF;
mem[16'hE7AE] = 8'h85;
mem[16'hE7AF] = 8'hA2;
mem[16'hE7B0] = 8'h45;
mem[16'hE7B1] = 8'hAA;
mem[16'hE7B2] = 8'h85;
mem[16'hE7B3] = 8'hAB;
mem[16'hE7B4] = 8'hA5;
mem[16'hE7B5] = 8'h9D;
mem[16'hE7B6] = 8'h4C;
mem[16'hE7B7] = 8'hC1;
mem[16'hE7B8] = 8'hE7;
mem[16'hE7B9] = 8'h20;
mem[16'hE7BA] = 8'hF0;
mem[16'hE7BB] = 8'hE8;
mem[16'hE7BC] = 8'h90;
mem[16'hE7BD] = 8'h3C;
mem[16'hE7BE] = 8'h20;
mem[16'hE7BF] = 8'hE3;
mem[16'hE7C0] = 8'hE9;
mem[16'hE7C1] = 8'hD0;
mem[16'hE7C2] = 8'h03;
mem[16'hE7C3] = 8'h4C;
mem[16'hE7C4] = 8'h53;
mem[16'hE7C5] = 8'hEB;
mem[16'hE7C6] = 8'hA6;
mem[16'hE7C7] = 8'hAC;
mem[16'hE7C8] = 8'h86;
mem[16'hE7C9] = 8'h92;
mem[16'hE7CA] = 8'hA2;
mem[16'hE7CB] = 8'hA5;
mem[16'hE7CC] = 8'hA5;
mem[16'hE7CD] = 8'hA5;
mem[16'hE7CE] = 8'hA8;
mem[16'hE7CF] = 8'hF0;
mem[16'hE7D0] = 8'hCE;
mem[16'hE7D1] = 8'h38;
mem[16'hE7D2] = 8'hE5;
mem[16'hE7D3] = 8'h9D;
mem[16'hE7D4] = 8'hF0;
mem[16'hE7D5] = 8'h24;
mem[16'hE7D6] = 8'h90;
mem[16'hE7D7] = 8'h12;
mem[16'hE7D8] = 8'h84;
mem[16'hE7D9] = 8'h9D;
mem[16'hE7DA] = 8'hA4;
mem[16'hE7DB] = 8'hAA;
mem[16'hE7DC] = 8'h84;
mem[16'hE7DD] = 8'hA2;
mem[16'hE7DE] = 8'h49;
mem[16'hE7DF] = 8'hFF;
mem[16'hE7E0] = 8'h69;
mem[16'hE7E1] = 8'h00;
mem[16'hE7E2] = 8'hA0;
mem[16'hE7E3] = 8'h00;
mem[16'hE7E4] = 8'h84;
mem[16'hE7E5] = 8'h92;
mem[16'hE7E6] = 8'hA2;
mem[16'hE7E7] = 8'h9D;
mem[16'hE7E8] = 8'hD0;
mem[16'hE7E9] = 8'h04;
mem[16'hE7EA] = 8'hA0;
mem[16'hE7EB] = 8'h00;
mem[16'hE7EC] = 8'h84;
mem[16'hE7ED] = 8'hAC;
mem[16'hE7EE] = 8'hC9;
mem[16'hE7EF] = 8'hF9;
mem[16'hE7F0] = 8'h30;
mem[16'hE7F1] = 8'hC7;
mem[16'hE7F2] = 8'hA8;
mem[16'hE7F3] = 8'hA5;
mem[16'hE7F4] = 8'hAC;
mem[16'hE7F5] = 8'h56;
mem[16'hE7F6] = 8'h01;
mem[16'hE7F7] = 8'h20;
mem[16'hE7F8] = 8'h07;
mem[16'hE7F9] = 8'hE9;
mem[16'hE7FA] = 8'h24;
mem[16'hE7FB] = 8'hAB;
mem[16'hE7FC] = 8'h10;
mem[16'hE7FD] = 8'h57;
mem[16'hE7FE] = 8'hA0;
mem[16'hE7FF] = 8'h9D;
mem[16'hE800] = 8'hE0;
mem[16'hE801] = 8'hA5;
mem[16'hE802] = 8'hF0;
mem[16'hE803] = 8'h02;
mem[16'hE804] = 8'hA0;
mem[16'hE805] = 8'hA5;
mem[16'hE806] = 8'h38;
mem[16'hE807] = 8'h49;
mem[16'hE808] = 8'hFF;
mem[16'hE809] = 8'h65;
mem[16'hE80A] = 8'h92;
mem[16'hE80B] = 8'h85;
mem[16'hE80C] = 8'hAC;
mem[16'hE80D] = 8'hB9;
mem[16'hE80E] = 8'h04;
mem[16'hE80F] = 8'h00;
mem[16'hE810] = 8'hF5;
mem[16'hE811] = 8'h04;
mem[16'hE812] = 8'h85;
mem[16'hE813] = 8'hA1;
mem[16'hE814] = 8'hB9;
mem[16'hE815] = 8'h03;
mem[16'hE816] = 8'h00;
mem[16'hE817] = 8'hF5;
mem[16'hE818] = 8'h03;
mem[16'hE819] = 8'h85;
mem[16'hE81A] = 8'hA0;
mem[16'hE81B] = 8'hB9;
mem[16'hE81C] = 8'h02;
mem[16'hE81D] = 8'h00;
mem[16'hE81E] = 8'hF5;
mem[16'hE81F] = 8'h02;
mem[16'hE820] = 8'h85;
mem[16'hE821] = 8'h9F;
mem[16'hE822] = 8'hB9;
mem[16'hE823] = 8'h01;
mem[16'hE824] = 8'h00;
mem[16'hE825] = 8'hF5;
mem[16'hE826] = 8'h01;
mem[16'hE827] = 8'h85;
mem[16'hE828] = 8'h9E;
mem[16'hE829] = 8'hB0;
mem[16'hE82A] = 8'h03;
mem[16'hE82B] = 8'h20;
mem[16'hE82C] = 8'h9E;
mem[16'hE82D] = 8'hE8;
mem[16'hE82E] = 8'hA0;
mem[16'hE82F] = 8'h00;
mem[16'hE830] = 8'h98;
mem[16'hE831] = 8'h18;
mem[16'hE832] = 8'hA6;
mem[16'hE833] = 8'h9E;
mem[16'hE834] = 8'hD0;
mem[16'hE835] = 8'h4A;
mem[16'hE836] = 8'hA6;
mem[16'hE837] = 8'h9F;
mem[16'hE838] = 8'h86;
mem[16'hE839] = 8'h9E;
mem[16'hE83A] = 8'hA6;
mem[16'hE83B] = 8'hA0;
mem[16'hE83C] = 8'h86;
mem[16'hE83D] = 8'h9F;
mem[16'hE83E] = 8'hA6;
mem[16'hE83F] = 8'hA1;
mem[16'hE840] = 8'h86;
mem[16'hE841] = 8'hA0;
mem[16'hE842] = 8'hA6;
mem[16'hE843] = 8'hAC;
mem[16'hE844] = 8'h86;
mem[16'hE845] = 8'hA1;
mem[16'hE846] = 8'h84;
mem[16'hE847] = 8'hAC;
mem[16'hE848] = 8'h69;
mem[16'hE849] = 8'h08;
mem[16'hE84A] = 8'hC9;
mem[16'hE84B] = 8'h20;
mem[16'hE84C] = 8'hD0;
mem[16'hE84D] = 8'hE4;
mem[16'hE84E] = 8'hA9;
mem[16'hE84F] = 8'h00;
mem[16'hE850] = 8'h85;
mem[16'hE851] = 8'h9D;
mem[16'hE852] = 8'h85;
mem[16'hE853] = 8'hA2;
mem[16'hE854] = 8'h60;
mem[16'hE855] = 8'h65;
mem[16'hE856] = 8'h92;
mem[16'hE857] = 8'h85;
mem[16'hE858] = 8'hAC;
mem[16'hE859] = 8'hA5;
mem[16'hE85A] = 8'hA1;
mem[16'hE85B] = 8'h65;
mem[16'hE85C] = 8'hA9;
mem[16'hE85D] = 8'h85;
mem[16'hE85E] = 8'hA1;
mem[16'hE85F] = 8'hA5;
mem[16'hE860] = 8'hA0;
mem[16'hE861] = 8'h65;
mem[16'hE862] = 8'hA8;
mem[16'hE863] = 8'h85;
mem[16'hE864] = 8'hA0;
mem[16'hE865] = 8'hA5;
mem[16'hE866] = 8'h9F;
mem[16'hE867] = 8'h65;
mem[16'hE868] = 8'hA7;
mem[16'hE869] = 8'h85;
mem[16'hE86A] = 8'h9F;
mem[16'hE86B] = 8'hA5;
mem[16'hE86C] = 8'h9E;
mem[16'hE86D] = 8'h65;
mem[16'hE86E] = 8'hA6;
mem[16'hE86F] = 8'h85;
mem[16'hE870] = 8'h9E;
mem[16'hE871] = 8'h4C;
mem[16'hE872] = 8'h8D;
mem[16'hE873] = 8'hE8;
mem[16'hE874] = 8'h69;
mem[16'hE875] = 8'h01;
mem[16'hE876] = 8'h06;
mem[16'hE877] = 8'hAC;
mem[16'hE878] = 8'h26;
mem[16'hE879] = 8'hA1;
mem[16'hE87A] = 8'h26;
mem[16'hE87B] = 8'hA0;
mem[16'hE87C] = 8'h26;
mem[16'hE87D] = 8'h9F;
mem[16'hE87E] = 8'h26;
mem[16'hE87F] = 8'h9E;
mem[16'hE880] = 8'h10;
mem[16'hE881] = 8'hF2;
mem[16'hE882] = 8'h38;
mem[16'hE883] = 8'hE5;
mem[16'hE884] = 8'h9D;
mem[16'hE885] = 8'hB0;
mem[16'hE886] = 8'hC7;
mem[16'hE887] = 8'h49;
mem[16'hE888] = 8'hFF;
mem[16'hE889] = 8'h69;
mem[16'hE88A] = 8'h01;
mem[16'hE88B] = 8'h85;
mem[16'hE88C] = 8'h9D;
mem[16'hE88D] = 8'h90;
mem[16'hE88E] = 8'h0E;
mem[16'hE88F] = 8'hE6;
mem[16'hE890] = 8'h9D;
mem[16'hE891] = 8'hF0;
mem[16'hE892] = 8'h42;
mem[16'hE893] = 8'h66;
mem[16'hE894] = 8'h9E;
mem[16'hE895] = 8'h66;
mem[16'hE896] = 8'h9F;
mem[16'hE897] = 8'h66;
mem[16'hE898] = 8'hA0;
mem[16'hE899] = 8'h66;
mem[16'hE89A] = 8'hA1;
mem[16'hE89B] = 8'h66;
mem[16'hE89C] = 8'hAC;
mem[16'hE89D] = 8'h60;
mem[16'hE89E] = 8'hA5;
mem[16'hE89F] = 8'hA2;
mem[16'hE8A0] = 8'h49;
mem[16'hE8A1] = 8'hFF;
mem[16'hE8A2] = 8'h85;
mem[16'hE8A3] = 8'hA2;
mem[16'hE8A4] = 8'hA5;
mem[16'hE8A5] = 8'h9E;
mem[16'hE8A6] = 8'h49;
mem[16'hE8A7] = 8'hFF;
mem[16'hE8A8] = 8'h85;
mem[16'hE8A9] = 8'h9E;
mem[16'hE8AA] = 8'hA5;
mem[16'hE8AB] = 8'h9F;
mem[16'hE8AC] = 8'h49;
mem[16'hE8AD] = 8'hFF;
mem[16'hE8AE] = 8'h85;
mem[16'hE8AF] = 8'h9F;
mem[16'hE8B0] = 8'hA5;
mem[16'hE8B1] = 8'hA0;
mem[16'hE8B2] = 8'h49;
mem[16'hE8B3] = 8'hFF;
mem[16'hE8B4] = 8'h85;
mem[16'hE8B5] = 8'hA0;
mem[16'hE8B6] = 8'hA5;
mem[16'hE8B7] = 8'hA1;
mem[16'hE8B8] = 8'h49;
mem[16'hE8B9] = 8'hFF;
mem[16'hE8BA] = 8'h85;
mem[16'hE8BB] = 8'hA1;
mem[16'hE8BC] = 8'hA5;
mem[16'hE8BD] = 8'hAC;
mem[16'hE8BE] = 8'h49;
mem[16'hE8BF] = 8'hFF;
mem[16'hE8C0] = 8'h85;
mem[16'hE8C1] = 8'hAC;
mem[16'hE8C2] = 8'hE6;
mem[16'hE8C3] = 8'hAC;
mem[16'hE8C4] = 8'hD0;
mem[16'hE8C5] = 8'h0E;
mem[16'hE8C6] = 8'hE6;
mem[16'hE8C7] = 8'hA1;
mem[16'hE8C8] = 8'hD0;
mem[16'hE8C9] = 8'h0A;
mem[16'hE8CA] = 8'hE6;
mem[16'hE8CB] = 8'hA0;
mem[16'hE8CC] = 8'hD0;
mem[16'hE8CD] = 8'h06;
mem[16'hE8CE] = 8'hE6;
mem[16'hE8CF] = 8'h9F;
mem[16'hE8D0] = 8'hD0;
mem[16'hE8D1] = 8'h02;
mem[16'hE8D2] = 8'hE6;
mem[16'hE8D3] = 8'h9E;
mem[16'hE8D4] = 8'h60;
mem[16'hE8D5] = 8'hA2;
mem[16'hE8D6] = 8'h45;
mem[16'hE8D7] = 8'h4C;
mem[16'hE8D8] = 8'h12;
mem[16'hE8D9] = 8'hD4;
mem[16'hE8DA] = 8'hA2;
mem[16'hE8DB] = 8'h61;
mem[16'hE8DC] = 8'hB4;
mem[16'hE8DD] = 8'h04;
mem[16'hE8DE] = 8'h84;
mem[16'hE8DF] = 8'hAC;
mem[16'hE8E0] = 8'hB4;
mem[16'hE8E1] = 8'h03;
mem[16'hE8E2] = 8'h94;
mem[16'hE8E3] = 8'h04;
mem[16'hE8E4] = 8'hB4;
mem[16'hE8E5] = 8'h02;
mem[16'hE8E6] = 8'h94;
mem[16'hE8E7] = 8'h03;
mem[16'hE8E8] = 8'hB4;
mem[16'hE8E9] = 8'h01;
mem[16'hE8EA] = 8'h94;
mem[16'hE8EB] = 8'h02;
mem[16'hE8EC] = 8'hA4;
mem[16'hE8ED] = 8'hA4;
mem[16'hE8EE] = 8'h94;
mem[16'hE8EF] = 8'h01;
mem[16'hE8F0] = 8'h69;
mem[16'hE8F1] = 8'h08;
mem[16'hE8F2] = 8'h30;
mem[16'hE8F3] = 8'hE8;
mem[16'hE8F4] = 8'hF0;
mem[16'hE8F5] = 8'hE6;
mem[16'hE8F6] = 8'hE9;
mem[16'hE8F7] = 8'h08;
mem[16'hE8F8] = 8'hA8;
mem[16'hE8F9] = 8'hA5;
mem[16'hE8FA] = 8'hAC;
mem[16'hE8FB] = 8'hB0;
mem[16'hE8FC] = 8'h14;
mem[16'hE8FD] = 8'h16;
mem[16'hE8FE] = 8'h01;
mem[16'hE8FF] = 8'h90;
mem[16'hE900] = 8'h02;
mem[16'hE901] = 8'hF6;
mem[16'hE902] = 8'h01;
mem[16'hE903] = 8'h76;
mem[16'hE904] = 8'h01;
mem[16'hE905] = 8'h76;
mem[16'hE906] = 8'h01;
mem[16'hE907] = 8'h76;
mem[16'hE908] = 8'h02;
mem[16'hE909] = 8'h76;
mem[16'hE90A] = 8'h03;
mem[16'hE90B] = 8'h76;
mem[16'hE90C] = 8'h04;
mem[16'hE90D] = 8'h6A;
mem[16'hE90E] = 8'hC8;
mem[16'hE90F] = 8'hD0;
mem[16'hE910] = 8'hEC;
mem[16'hE911] = 8'h18;
mem[16'hE912] = 8'h60;
mem[16'hE913] = 8'h81;
mem[16'hE914] = 8'h00;
mem[16'hE915] = 8'h00;
mem[16'hE916] = 8'h00;
mem[16'hE917] = 8'h00;
mem[16'hE918] = 8'h03;
mem[16'hE919] = 8'h7F;
mem[16'hE91A] = 8'h5E;
mem[16'hE91B] = 8'h56;
mem[16'hE91C] = 8'hCB;
mem[16'hE91D] = 8'h79;
mem[16'hE91E] = 8'h80;
mem[16'hE91F] = 8'h13;
mem[16'hE920] = 8'h9B;
mem[16'hE921] = 8'h0B;
mem[16'hE922] = 8'h64;
mem[16'hE923] = 8'h80;
mem[16'hE924] = 8'h76;
mem[16'hE925] = 8'h38;
mem[16'hE926] = 8'h93;
mem[16'hE927] = 8'h16;
mem[16'hE928] = 8'h82;
mem[16'hE929] = 8'h38;
mem[16'hE92A] = 8'hAA;
mem[16'hE92B] = 8'h3B;
mem[16'hE92C] = 8'h20;
mem[16'hE92D] = 8'h80;
mem[16'hE92E] = 8'h35;
mem[16'hE92F] = 8'h04;
mem[16'hE930] = 8'hF3;
mem[16'hE931] = 8'h34;
mem[16'hE932] = 8'h81;
mem[16'hE933] = 8'h35;
mem[16'hE934] = 8'h04;
mem[16'hE935] = 8'hF3;
mem[16'hE936] = 8'h34;
mem[16'hE937] = 8'h80;
mem[16'hE938] = 8'h80;
mem[16'hE939] = 8'h00;
mem[16'hE93A] = 8'h00;
mem[16'hE93B] = 8'h00;
mem[16'hE93C] = 8'h80;
mem[16'hE93D] = 8'h31;
mem[16'hE93E] = 8'h72;
mem[16'hE93F] = 8'h17;
mem[16'hE940] = 8'hF8;
mem[16'hE941] = 8'h20;
mem[16'hE942] = 8'h82;
mem[16'hE943] = 8'hEB;
mem[16'hE944] = 8'hF0;
mem[16'hE945] = 8'h02;
mem[16'hE946] = 8'h10;
mem[16'hE947] = 8'h03;
mem[16'hE948] = 8'h4C;
mem[16'hE949] = 8'h99;
mem[16'hE94A] = 8'hE1;
mem[16'hE94B] = 8'hA5;
mem[16'hE94C] = 8'h9D;
mem[16'hE94D] = 8'hE9;
mem[16'hE94E] = 8'h7F;
mem[16'hE94F] = 8'h48;
mem[16'hE950] = 8'hA9;
mem[16'hE951] = 8'h80;
mem[16'hE952] = 8'h85;
mem[16'hE953] = 8'h9D;
mem[16'hE954] = 8'hA9;
mem[16'hE955] = 8'h2D;
mem[16'hE956] = 8'hA0;
mem[16'hE957] = 8'hE9;
mem[16'hE958] = 8'h20;
mem[16'hE959] = 8'hBE;
mem[16'hE95A] = 8'hE7;
mem[16'hE95B] = 8'hA9;
mem[16'hE95C] = 8'h32;
mem[16'hE95D] = 8'hA0;
mem[16'hE95E] = 8'hE9;
mem[16'hE95F] = 8'h20;
mem[16'hE960] = 8'h66;
mem[16'hE961] = 8'hEA;
mem[16'hE962] = 8'hA9;
mem[16'hE963] = 8'h13;
mem[16'hE964] = 8'hA0;
mem[16'hE965] = 8'hE9;
mem[16'hE966] = 8'h20;
mem[16'hE967] = 8'hA7;
mem[16'hE968] = 8'hE7;
mem[16'hE969] = 8'hA9;
mem[16'hE96A] = 8'h18;
mem[16'hE96B] = 8'hA0;
mem[16'hE96C] = 8'hE9;
mem[16'hE96D] = 8'h20;
mem[16'hE96E] = 8'h5C;
mem[16'hE96F] = 8'hEF;
mem[16'hE970] = 8'hA9;
mem[16'hE971] = 8'h37;
mem[16'hE972] = 8'hA0;
mem[16'hE973] = 8'hE9;
mem[16'hE974] = 8'h20;
mem[16'hE975] = 8'hBE;
mem[16'hE976] = 8'hE7;
mem[16'hE977] = 8'h68;
mem[16'hE978] = 8'h20;
mem[16'hE979] = 8'hD5;
mem[16'hE97A] = 8'hEC;
mem[16'hE97B] = 8'hA9;
mem[16'hE97C] = 8'h3C;
mem[16'hE97D] = 8'hA0;
mem[16'hE97E] = 8'hE9;
mem[16'hE97F] = 8'h20;
mem[16'hE980] = 8'hE3;
mem[16'hE981] = 8'hE9;
mem[16'hE982] = 8'hD0;
mem[16'hE983] = 8'h03;
mem[16'hE984] = 8'h4C;
mem[16'hE985] = 8'hE2;
mem[16'hE986] = 8'hE9;
mem[16'hE987] = 8'h20;
mem[16'hE988] = 8'h0E;
mem[16'hE989] = 8'hEA;
mem[16'hE98A] = 8'hA9;
mem[16'hE98B] = 8'h00;
mem[16'hE98C] = 8'h85;
mem[16'hE98D] = 8'h62;
mem[16'hE98E] = 8'h85;
mem[16'hE98F] = 8'h63;
mem[16'hE990] = 8'h85;
mem[16'hE991] = 8'h64;
mem[16'hE992] = 8'h85;
mem[16'hE993] = 8'h65;
mem[16'hE994] = 8'hA5;
mem[16'hE995] = 8'hAC;
mem[16'hE996] = 8'h20;
mem[16'hE997] = 8'hB0;
mem[16'hE998] = 8'hE9;
mem[16'hE999] = 8'hA5;
mem[16'hE99A] = 8'hA1;
mem[16'hE99B] = 8'h20;
mem[16'hE99C] = 8'hB0;
mem[16'hE99D] = 8'hE9;
mem[16'hE99E] = 8'hA5;
mem[16'hE99F] = 8'hA0;
mem[16'hE9A0] = 8'h20;
mem[16'hE9A1] = 8'hB0;
mem[16'hE9A2] = 8'hE9;
mem[16'hE9A3] = 8'hA5;
mem[16'hE9A4] = 8'h9F;
mem[16'hE9A5] = 8'h20;
mem[16'hE9A6] = 8'hB0;
mem[16'hE9A7] = 8'hE9;
mem[16'hE9A8] = 8'hA5;
mem[16'hE9A9] = 8'h9E;
mem[16'hE9AA] = 8'h20;
mem[16'hE9AB] = 8'hB5;
mem[16'hE9AC] = 8'hE9;
mem[16'hE9AD] = 8'h4C;
mem[16'hE9AE] = 8'hE6;
mem[16'hE9AF] = 8'hEA;
mem[16'hE9B0] = 8'hD0;
mem[16'hE9B1] = 8'h03;
mem[16'hE9B2] = 8'h4C;
mem[16'hE9B3] = 8'hDA;
mem[16'hE9B4] = 8'hE8;
mem[16'hE9B5] = 8'h4A;
mem[16'hE9B6] = 8'h09;
mem[16'hE9B7] = 8'h80;
mem[16'hE9B8] = 8'hA8;
mem[16'hE9B9] = 8'h90;
mem[16'hE9BA] = 8'h19;
mem[16'hE9BB] = 8'h18;
mem[16'hE9BC] = 8'hA5;
mem[16'hE9BD] = 8'h65;
mem[16'hE9BE] = 8'h65;
mem[16'hE9BF] = 8'hA9;
mem[16'hE9C0] = 8'h85;
mem[16'hE9C1] = 8'h65;
mem[16'hE9C2] = 8'hA5;
mem[16'hE9C3] = 8'h64;
mem[16'hE9C4] = 8'h65;
mem[16'hE9C5] = 8'hA8;
mem[16'hE9C6] = 8'h85;
mem[16'hE9C7] = 8'h64;
mem[16'hE9C8] = 8'hA5;
mem[16'hE9C9] = 8'h63;
mem[16'hE9CA] = 8'h65;
mem[16'hE9CB] = 8'hA7;
mem[16'hE9CC] = 8'h85;
mem[16'hE9CD] = 8'h63;
mem[16'hE9CE] = 8'hA5;
mem[16'hE9CF] = 8'h62;
mem[16'hE9D0] = 8'h65;
mem[16'hE9D1] = 8'hA6;
mem[16'hE9D2] = 8'h85;
mem[16'hE9D3] = 8'h62;
mem[16'hE9D4] = 8'h66;
mem[16'hE9D5] = 8'h62;
mem[16'hE9D6] = 8'h66;
mem[16'hE9D7] = 8'h63;
mem[16'hE9D8] = 8'h66;
mem[16'hE9D9] = 8'h64;
mem[16'hE9DA] = 8'h66;
mem[16'hE9DB] = 8'h65;
mem[16'hE9DC] = 8'h66;
mem[16'hE9DD] = 8'hAC;
mem[16'hE9DE] = 8'h98;
mem[16'hE9DF] = 8'h4A;
mem[16'hE9E0] = 8'hD0;
mem[16'hE9E1] = 8'hD6;
mem[16'hE9E2] = 8'h60;
mem[16'hE9E3] = 8'h85;
mem[16'hE9E4] = 8'h5E;
mem[16'hE9E5] = 8'h84;
mem[16'hE9E6] = 8'h5F;
mem[16'hE9E7] = 8'hA0;
mem[16'hE9E8] = 8'h04;
mem[16'hE9E9] = 8'hB1;
mem[16'hE9EA] = 8'h5E;
mem[16'hE9EB] = 8'h85;
mem[16'hE9EC] = 8'hA9;
mem[16'hE9ED] = 8'h88;
mem[16'hE9EE] = 8'hB1;
mem[16'hE9EF] = 8'h5E;
mem[16'hE9F0] = 8'h85;
mem[16'hE9F1] = 8'hA8;
mem[16'hE9F2] = 8'h88;
mem[16'hE9F3] = 8'hB1;
mem[16'hE9F4] = 8'h5E;
mem[16'hE9F5] = 8'h85;
mem[16'hE9F6] = 8'hA7;
mem[16'hE9F7] = 8'h88;
mem[16'hE9F8] = 8'hB1;
mem[16'hE9F9] = 8'h5E;
mem[16'hE9FA] = 8'h85;
mem[16'hE9FB] = 8'hAA;
mem[16'hE9FC] = 8'h45;
mem[16'hE9FD] = 8'hA2;
mem[16'hE9FE] = 8'h85;
mem[16'hE9FF] = 8'hAB;
mem[16'hEA00] = 8'hA5;
mem[16'hEA01] = 8'hAA;
mem[16'hEA02] = 8'h09;
mem[16'hEA03] = 8'h80;
mem[16'hEA04] = 8'h85;
mem[16'hEA05] = 8'hA6;
mem[16'hEA06] = 8'h88;
mem[16'hEA07] = 8'hB1;
mem[16'hEA08] = 8'h5E;
mem[16'hEA09] = 8'h85;
mem[16'hEA0A] = 8'hA5;
mem[16'hEA0B] = 8'hA5;
mem[16'hEA0C] = 8'h9D;
mem[16'hEA0D] = 8'h60;
mem[16'hEA0E] = 8'hA5;
mem[16'hEA0F] = 8'hA5;
mem[16'hEA10] = 8'hF0;
mem[16'hEA11] = 8'h1F;
mem[16'hEA12] = 8'h18;
mem[16'hEA13] = 8'h65;
mem[16'hEA14] = 8'h9D;
mem[16'hEA15] = 8'h90;
mem[16'hEA16] = 8'h04;
mem[16'hEA17] = 8'h30;
mem[16'hEA18] = 8'h1D;
mem[16'hEA19] = 8'h18;
mem[16'hEA1A] = 8'h2C;
mem[16'hEA1B] = 8'h10;
mem[16'hEA1C] = 8'h14;
mem[16'hEA1D] = 8'h69;
mem[16'hEA1E] = 8'h80;
mem[16'hEA1F] = 8'h85;
mem[16'hEA20] = 8'h9D;
mem[16'hEA21] = 8'hD0;
mem[16'hEA22] = 8'h03;
mem[16'hEA23] = 8'h4C;
mem[16'hEA24] = 8'h52;
mem[16'hEA25] = 8'hE8;
mem[16'hEA26] = 8'hA5;
mem[16'hEA27] = 8'hAB;
mem[16'hEA28] = 8'h85;
mem[16'hEA29] = 8'hA2;
mem[16'hEA2A] = 8'h60;
mem[16'hEA2B] = 8'hA5;
mem[16'hEA2C] = 8'hA2;
mem[16'hEA2D] = 8'h49;
mem[16'hEA2E] = 8'hFF;
mem[16'hEA2F] = 8'h30;
mem[16'hEA30] = 8'h05;
mem[16'hEA31] = 8'h68;
mem[16'hEA32] = 8'h68;
mem[16'hEA33] = 8'h4C;
mem[16'hEA34] = 8'h4E;
mem[16'hEA35] = 8'hE8;
mem[16'hEA36] = 8'h4C;
mem[16'hEA37] = 8'hD5;
mem[16'hEA38] = 8'hE8;
mem[16'hEA39] = 8'h20;
mem[16'hEA3A] = 8'h63;
mem[16'hEA3B] = 8'hEB;
mem[16'hEA3C] = 8'hAA;
mem[16'hEA3D] = 8'hF0;
mem[16'hEA3E] = 8'h10;
mem[16'hEA3F] = 8'h18;
mem[16'hEA40] = 8'h69;
mem[16'hEA41] = 8'h02;
mem[16'hEA42] = 8'hB0;
mem[16'hEA43] = 8'hF2;
mem[16'hEA44] = 8'hA2;
mem[16'hEA45] = 8'h00;
mem[16'hEA46] = 8'h86;
mem[16'hEA47] = 8'hAB;
mem[16'hEA48] = 8'h20;
mem[16'hEA49] = 8'hCE;
mem[16'hEA4A] = 8'hE7;
mem[16'hEA4B] = 8'hE6;
mem[16'hEA4C] = 8'h9D;
mem[16'hEA4D] = 8'hF0;
mem[16'hEA4E] = 8'hE7;
mem[16'hEA4F] = 8'h60;
mem[16'hEA50] = 8'h84;
mem[16'hEA51] = 8'h20;
mem[16'hEA52] = 8'h00;
mem[16'hEA53] = 8'h00;
mem[16'hEA54] = 8'h00;
mem[16'hEA55] = 8'h20;
mem[16'hEA56] = 8'h63;
mem[16'hEA57] = 8'hEB;
mem[16'hEA58] = 8'hA9;
mem[16'hEA59] = 8'h50;
mem[16'hEA5A] = 8'hA0;
mem[16'hEA5B] = 8'hEA;
mem[16'hEA5C] = 8'hA2;
mem[16'hEA5D] = 8'h00;
mem[16'hEA5E] = 8'h86;
mem[16'hEA5F] = 8'hAB;
mem[16'hEA60] = 8'h20;
mem[16'hEA61] = 8'hF9;
mem[16'hEA62] = 8'hEA;
mem[16'hEA63] = 8'h4C;
mem[16'hEA64] = 8'h69;
mem[16'hEA65] = 8'hEA;
mem[16'hEA66] = 8'h20;
mem[16'hEA67] = 8'hE3;
mem[16'hEA68] = 8'hE9;
mem[16'hEA69] = 8'hF0;
mem[16'hEA6A] = 8'h76;
mem[16'hEA6B] = 8'h20;
mem[16'hEA6C] = 8'h72;
mem[16'hEA6D] = 8'hEB;
mem[16'hEA6E] = 8'hA9;
mem[16'hEA6F] = 8'h00;
mem[16'hEA70] = 8'h38;
mem[16'hEA71] = 8'hE5;
mem[16'hEA72] = 8'h9D;
mem[16'hEA73] = 8'h85;
mem[16'hEA74] = 8'h9D;
mem[16'hEA75] = 8'h20;
mem[16'hEA76] = 8'h0E;
mem[16'hEA77] = 8'hEA;
mem[16'hEA78] = 8'hE6;
mem[16'hEA79] = 8'h9D;
mem[16'hEA7A] = 8'hF0;
mem[16'hEA7B] = 8'hBA;
mem[16'hEA7C] = 8'hA2;
mem[16'hEA7D] = 8'hFC;
mem[16'hEA7E] = 8'hA9;
mem[16'hEA7F] = 8'h01;
mem[16'hEA80] = 8'hA4;
mem[16'hEA81] = 8'hA6;
mem[16'hEA82] = 8'hC4;
mem[16'hEA83] = 8'h9E;
mem[16'hEA84] = 8'hD0;
mem[16'hEA85] = 8'h10;
mem[16'hEA86] = 8'hA4;
mem[16'hEA87] = 8'hA7;
mem[16'hEA88] = 8'hC4;
mem[16'hEA89] = 8'h9F;
mem[16'hEA8A] = 8'hD0;
mem[16'hEA8B] = 8'h0A;
mem[16'hEA8C] = 8'hA4;
mem[16'hEA8D] = 8'hA8;
mem[16'hEA8E] = 8'hC4;
mem[16'hEA8F] = 8'hA0;
mem[16'hEA90] = 8'hD0;
mem[16'hEA91] = 8'h04;
mem[16'hEA92] = 8'hA4;
mem[16'hEA93] = 8'hA9;
mem[16'hEA94] = 8'hC4;
mem[16'hEA95] = 8'hA1;
mem[16'hEA96] = 8'h08;
mem[16'hEA97] = 8'h2A;
mem[16'hEA98] = 8'h90;
mem[16'hEA99] = 8'h09;
mem[16'hEA9A] = 8'hE8;
mem[16'hEA9B] = 8'h95;
mem[16'hEA9C] = 8'h65;
mem[16'hEA9D] = 8'hF0;
mem[16'hEA9E] = 8'h32;
mem[16'hEA9F] = 8'h10;
mem[16'hEAA0] = 8'h34;
mem[16'hEAA1] = 8'hA9;
mem[16'hEAA2] = 8'h01;
mem[16'hEAA3] = 8'h28;
mem[16'hEAA4] = 8'hB0;
mem[16'hEAA5] = 8'h0E;
mem[16'hEAA6] = 8'h06;
mem[16'hEAA7] = 8'hA9;
mem[16'hEAA8] = 8'h26;
mem[16'hEAA9] = 8'hA8;
mem[16'hEAAA] = 8'h26;
mem[16'hEAAB] = 8'hA7;
mem[16'hEAAC] = 8'h26;
mem[16'hEAAD] = 8'hA6;
mem[16'hEAAE] = 8'hB0;
mem[16'hEAAF] = 8'hE6;
mem[16'hEAB0] = 8'h30;
mem[16'hEAB1] = 8'hCE;
mem[16'hEAB2] = 8'h10;
mem[16'hEAB3] = 8'hE2;
mem[16'hEAB4] = 8'hA8;
mem[16'hEAB5] = 8'hA5;
mem[16'hEAB6] = 8'hA9;
mem[16'hEAB7] = 8'hE5;
mem[16'hEAB8] = 8'hA1;
mem[16'hEAB9] = 8'h85;
mem[16'hEABA] = 8'hA9;
mem[16'hEABB] = 8'hA5;
mem[16'hEABC] = 8'hA8;
mem[16'hEABD] = 8'hE5;
mem[16'hEABE] = 8'hA0;
mem[16'hEABF] = 8'h85;
mem[16'hEAC0] = 8'hA8;
mem[16'hEAC1] = 8'hA5;
mem[16'hEAC2] = 8'hA7;
mem[16'hEAC3] = 8'hE5;
mem[16'hEAC4] = 8'h9F;
mem[16'hEAC5] = 8'h85;
mem[16'hEAC6] = 8'hA7;
mem[16'hEAC7] = 8'hA5;
mem[16'hEAC8] = 8'hA6;
mem[16'hEAC9] = 8'hE5;
mem[16'hEACA] = 8'h9E;
mem[16'hEACB] = 8'h85;
mem[16'hEACC] = 8'hA6;
mem[16'hEACD] = 8'h98;
mem[16'hEACE] = 8'h4C;
mem[16'hEACF] = 8'hA6;
mem[16'hEAD0] = 8'hEA;
mem[16'hEAD1] = 8'hA9;
mem[16'hEAD2] = 8'h40;
mem[16'hEAD3] = 8'hD0;
mem[16'hEAD4] = 8'hCE;
mem[16'hEAD5] = 8'h0A;
mem[16'hEAD6] = 8'h0A;
mem[16'hEAD7] = 8'h0A;
mem[16'hEAD8] = 8'h0A;
mem[16'hEAD9] = 8'h0A;
mem[16'hEADA] = 8'h0A;
mem[16'hEADB] = 8'h85;
mem[16'hEADC] = 8'hAC;
mem[16'hEADD] = 8'h28;
mem[16'hEADE] = 8'h4C;
mem[16'hEADF] = 8'hE6;
mem[16'hEAE0] = 8'hEA;
mem[16'hEAE1] = 8'hA2;
mem[16'hEAE2] = 8'h85;
mem[16'hEAE3] = 8'h4C;
mem[16'hEAE4] = 8'h12;
mem[16'hEAE5] = 8'hD4;
mem[16'hEAE6] = 8'hA5;
mem[16'hEAE7] = 8'h62;
mem[16'hEAE8] = 8'h85;
mem[16'hEAE9] = 8'h9E;
mem[16'hEAEA] = 8'hA5;
mem[16'hEAEB] = 8'h63;
mem[16'hEAEC] = 8'h85;
mem[16'hEAED] = 8'h9F;
mem[16'hEAEE] = 8'hA5;
mem[16'hEAEF] = 8'h64;
mem[16'hEAF0] = 8'h85;
mem[16'hEAF1] = 8'hA0;
mem[16'hEAF2] = 8'hA5;
mem[16'hEAF3] = 8'h65;
mem[16'hEAF4] = 8'h85;
mem[16'hEAF5] = 8'hA1;
mem[16'hEAF6] = 8'h4C;
mem[16'hEAF7] = 8'h2E;
mem[16'hEAF8] = 8'hE8;
mem[16'hEAF9] = 8'h85;
mem[16'hEAFA] = 8'h5E;
mem[16'hEAFB] = 8'h84;
mem[16'hEAFC] = 8'h5F;
mem[16'hEAFD] = 8'hA0;
mem[16'hEAFE] = 8'h04;
mem[16'hEAFF] = 8'hB1;
mem[16'hEB00] = 8'h5E;
mem[16'hEB01] = 8'h85;
mem[16'hEB02] = 8'hA1;
mem[16'hEB03] = 8'h88;
mem[16'hEB04] = 8'hB1;
mem[16'hEB05] = 8'h5E;
mem[16'hEB06] = 8'h85;
mem[16'hEB07] = 8'hA0;
mem[16'hEB08] = 8'h88;
mem[16'hEB09] = 8'hB1;
mem[16'hEB0A] = 8'h5E;
mem[16'hEB0B] = 8'h85;
mem[16'hEB0C] = 8'h9F;
mem[16'hEB0D] = 8'h88;
mem[16'hEB0E] = 8'hB1;
mem[16'hEB0F] = 8'h5E;
mem[16'hEB10] = 8'h85;
mem[16'hEB11] = 8'hA2;
mem[16'hEB12] = 8'h09;
mem[16'hEB13] = 8'h80;
mem[16'hEB14] = 8'h85;
mem[16'hEB15] = 8'h9E;
mem[16'hEB16] = 8'h88;
mem[16'hEB17] = 8'hB1;
mem[16'hEB18] = 8'h5E;
mem[16'hEB19] = 8'h85;
mem[16'hEB1A] = 8'h9D;
mem[16'hEB1B] = 8'h84;
mem[16'hEB1C] = 8'hAC;
mem[16'hEB1D] = 8'h60;
mem[16'hEB1E] = 8'hA2;
mem[16'hEB1F] = 8'h98;
mem[16'hEB20] = 8'h2C;
mem[16'hEB21] = 8'hA2;
mem[16'hEB22] = 8'h93;
mem[16'hEB23] = 8'hA0;
mem[16'hEB24] = 8'h00;
mem[16'hEB25] = 8'hF0;
mem[16'hEB26] = 8'h04;
mem[16'hEB27] = 8'hA6;
mem[16'hEB28] = 8'h85;
mem[16'hEB29] = 8'hA4;
mem[16'hEB2A] = 8'h86;
mem[16'hEB2B] = 8'h20;
mem[16'hEB2C] = 8'h72;
mem[16'hEB2D] = 8'hEB;
mem[16'hEB2E] = 8'h86;
mem[16'hEB2F] = 8'h5E;
mem[16'hEB30] = 8'h84;
mem[16'hEB31] = 8'h5F;
mem[16'hEB32] = 8'hA0;
mem[16'hEB33] = 8'h04;
mem[16'hEB34] = 8'hA5;
mem[16'hEB35] = 8'hA1;
mem[16'hEB36] = 8'h91;
mem[16'hEB37] = 8'h5E;
mem[16'hEB38] = 8'h88;
mem[16'hEB39] = 8'hA5;
mem[16'hEB3A] = 8'hA0;
mem[16'hEB3B] = 8'h91;
mem[16'hEB3C] = 8'h5E;
mem[16'hEB3D] = 8'h88;
mem[16'hEB3E] = 8'hA5;
mem[16'hEB3F] = 8'h9F;
mem[16'hEB40] = 8'h91;
mem[16'hEB41] = 8'h5E;
mem[16'hEB42] = 8'h88;
mem[16'hEB43] = 8'hA5;
mem[16'hEB44] = 8'hA2;
mem[16'hEB45] = 8'h09;
mem[16'hEB46] = 8'h7F;
mem[16'hEB47] = 8'h25;
mem[16'hEB48] = 8'h9E;
mem[16'hEB49] = 8'h91;
mem[16'hEB4A] = 8'h5E;
mem[16'hEB4B] = 8'h88;
mem[16'hEB4C] = 8'hA5;
mem[16'hEB4D] = 8'h9D;
mem[16'hEB4E] = 8'h91;
mem[16'hEB4F] = 8'h5E;
mem[16'hEB50] = 8'h84;
mem[16'hEB51] = 8'hAC;
mem[16'hEB52] = 8'h60;
mem[16'hEB53] = 8'hA5;
mem[16'hEB54] = 8'hAA;
mem[16'hEB55] = 8'h85;
mem[16'hEB56] = 8'hA2;
mem[16'hEB57] = 8'hA2;
mem[16'hEB58] = 8'h05;
mem[16'hEB59] = 8'hB5;
mem[16'hEB5A] = 8'hA4;
mem[16'hEB5B] = 8'h95;
mem[16'hEB5C] = 8'h9C;
mem[16'hEB5D] = 8'hCA;
mem[16'hEB5E] = 8'hD0;
mem[16'hEB5F] = 8'hF9;
mem[16'hEB60] = 8'h86;
mem[16'hEB61] = 8'hAC;
mem[16'hEB62] = 8'h60;
mem[16'hEB63] = 8'h20;
mem[16'hEB64] = 8'h72;
mem[16'hEB65] = 8'hEB;
mem[16'hEB66] = 8'hA2;
mem[16'hEB67] = 8'h06;
mem[16'hEB68] = 8'hB5;
mem[16'hEB69] = 8'h9C;
mem[16'hEB6A] = 8'h95;
mem[16'hEB6B] = 8'hA4;
mem[16'hEB6C] = 8'hCA;
mem[16'hEB6D] = 8'hD0;
mem[16'hEB6E] = 8'hF9;
mem[16'hEB6F] = 8'h86;
mem[16'hEB70] = 8'hAC;
mem[16'hEB71] = 8'h60;
mem[16'hEB72] = 8'hA5;
mem[16'hEB73] = 8'h9D;
mem[16'hEB74] = 8'hF0;
mem[16'hEB75] = 8'hFB;
mem[16'hEB76] = 8'h06;
mem[16'hEB77] = 8'hAC;
mem[16'hEB78] = 8'h90;
mem[16'hEB79] = 8'hF7;
mem[16'hEB7A] = 8'h20;
mem[16'hEB7B] = 8'hC6;
mem[16'hEB7C] = 8'hE8;
mem[16'hEB7D] = 8'hD0;
mem[16'hEB7E] = 8'hF2;
mem[16'hEB7F] = 8'h4C;
mem[16'hEB80] = 8'h8F;
mem[16'hEB81] = 8'hE8;
mem[16'hEB82] = 8'hA5;
mem[16'hEB83] = 8'h9D;
mem[16'hEB84] = 8'hF0;
mem[16'hEB85] = 8'h09;
mem[16'hEB86] = 8'hA5;
mem[16'hEB87] = 8'hA2;
mem[16'hEB88] = 8'h2A;
mem[16'hEB89] = 8'hA9;
mem[16'hEB8A] = 8'hFF;
mem[16'hEB8B] = 8'hB0;
mem[16'hEB8C] = 8'h02;
mem[16'hEB8D] = 8'hA9;
mem[16'hEB8E] = 8'h01;
mem[16'hEB8F] = 8'h60;
mem[16'hEB90] = 8'h20;
mem[16'hEB91] = 8'h82;
mem[16'hEB92] = 8'hEB;
mem[16'hEB93] = 8'h85;
mem[16'hEB94] = 8'h9E;
mem[16'hEB95] = 8'hA9;
mem[16'hEB96] = 8'h00;
mem[16'hEB97] = 8'h85;
mem[16'hEB98] = 8'h9F;
mem[16'hEB99] = 8'hA2;
mem[16'hEB9A] = 8'h88;
mem[16'hEB9B] = 8'hA5;
mem[16'hEB9C] = 8'h9E;
mem[16'hEB9D] = 8'h49;
mem[16'hEB9E] = 8'hFF;
mem[16'hEB9F] = 8'h2A;
mem[16'hEBA0] = 8'hA9;
mem[16'hEBA1] = 8'h00;
mem[16'hEBA2] = 8'h85;
mem[16'hEBA3] = 8'hA1;
mem[16'hEBA4] = 8'h85;
mem[16'hEBA5] = 8'hA0;
mem[16'hEBA6] = 8'h86;
mem[16'hEBA7] = 8'h9D;
mem[16'hEBA8] = 8'h85;
mem[16'hEBA9] = 8'hAC;
mem[16'hEBAA] = 8'h85;
mem[16'hEBAB] = 8'hA2;
mem[16'hEBAC] = 8'h4C;
mem[16'hEBAD] = 8'h29;
mem[16'hEBAE] = 8'hE8;
mem[16'hEBAF] = 8'h46;
mem[16'hEBB0] = 8'hA2;
mem[16'hEBB1] = 8'h60;
mem[16'hEBB2] = 8'h85;
mem[16'hEBB3] = 8'h60;
mem[16'hEBB4] = 8'h84;
mem[16'hEBB5] = 8'h61;
mem[16'hEBB6] = 8'hA0;
mem[16'hEBB7] = 8'h00;
mem[16'hEBB8] = 8'hB1;
mem[16'hEBB9] = 8'h60;
mem[16'hEBBA] = 8'hC8;
mem[16'hEBBB] = 8'hAA;
mem[16'hEBBC] = 8'hF0;
mem[16'hEBBD] = 8'hC4;
mem[16'hEBBE] = 8'hB1;
mem[16'hEBBF] = 8'h60;
mem[16'hEBC0] = 8'h45;
mem[16'hEBC1] = 8'hA2;
mem[16'hEBC2] = 8'h30;
mem[16'hEBC3] = 8'hC2;
mem[16'hEBC4] = 8'hE4;
mem[16'hEBC5] = 8'h9D;
mem[16'hEBC6] = 8'hD0;
mem[16'hEBC7] = 8'h21;
mem[16'hEBC8] = 8'hB1;
mem[16'hEBC9] = 8'h60;
mem[16'hEBCA] = 8'h09;
mem[16'hEBCB] = 8'h80;
mem[16'hEBCC] = 8'hC5;
mem[16'hEBCD] = 8'h9E;
mem[16'hEBCE] = 8'hD0;
mem[16'hEBCF] = 8'h19;
mem[16'hEBD0] = 8'hC8;
mem[16'hEBD1] = 8'hB1;
mem[16'hEBD2] = 8'h60;
mem[16'hEBD3] = 8'hC5;
mem[16'hEBD4] = 8'h9F;
mem[16'hEBD5] = 8'hD0;
mem[16'hEBD6] = 8'h12;
mem[16'hEBD7] = 8'hC8;
mem[16'hEBD8] = 8'hB1;
mem[16'hEBD9] = 8'h60;
mem[16'hEBDA] = 8'hC5;
mem[16'hEBDB] = 8'hA0;
mem[16'hEBDC] = 8'hD0;
mem[16'hEBDD] = 8'h0B;
mem[16'hEBDE] = 8'hC8;
mem[16'hEBDF] = 8'hA9;
mem[16'hEBE0] = 8'h7F;
mem[16'hEBE1] = 8'hC5;
mem[16'hEBE2] = 8'hAC;
mem[16'hEBE3] = 8'hB1;
mem[16'hEBE4] = 8'h60;
mem[16'hEBE5] = 8'hE5;
mem[16'hEBE6] = 8'hA1;
mem[16'hEBE7] = 8'hF0;
mem[16'hEBE8] = 8'h28;
mem[16'hEBE9] = 8'hA5;
mem[16'hEBEA] = 8'hA2;
mem[16'hEBEB] = 8'h90;
mem[16'hEBEC] = 8'h02;
mem[16'hEBED] = 8'h49;
mem[16'hEBEE] = 8'hFF;
mem[16'hEBEF] = 8'h4C;
mem[16'hEBF0] = 8'h88;
mem[16'hEBF1] = 8'hEB;
mem[16'hEBF2] = 8'hA5;
mem[16'hEBF3] = 8'h9D;
mem[16'hEBF4] = 8'hF0;
mem[16'hEBF5] = 8'h4A;
mem[16'hEBF6] = 8'h38;
mem[16'hEBF7] = 8'hE9;
mem[16'hEBF8] = 8'hA0;
mem[16'hEBF9] = 8'h24;
mem[16'hEBFA] = 8'hA2;
mem[16'hEBFB] = 8'h10;
mem[16'hEBFC] = 8'h09;
mem[16'hEBFD] = 8'hAA;
mem[16'hEBFE] = 8'hA9;
mem[16'hEBFF] = 8'hFF;
mem[16'hEC00] = 8'h85;
mem[16'hEC01] = 8'hA4;
mem[16'hEC02] = 8'h20;
mem[16'hEC03] = 8'hA4;
mem[16'hEC04] = 8'hE8;
mem[16'hEC05] = 8'h8A;
mem[16'hEC06] = 8'hA2;
mem[16'hEC07] = 8'h9D;
mem[16'hEC08] = 8'hC9;
mem[16'hEC09] = 8'hF9;
mem[16'hEC0A] = 8'h10;
mem[16'hEC0B] = 8'h06;
mem[16'hEC0C] = 8'h20;
mem[16'hEC0D] = 8'hF0;
mem[16'hEC0E] = 8'hE8;
mem[16'hEC0F] = 8'h84;
mem[16'hEC10] = 8'hA4;
mem[16'hEC11] = 8'h60;
mem[16'hEC12] = 8'hA8;
mem[16'hEC13] = 8'hA5;
mem[16'hEC14] = 8'hA2;
mem[16'hEC15] = 8'h29;
mem[16'hEC16] = 8'h80;
mem[16'hEC17] = 8'h46;
mem[16'hEC18] = 8'h9E;
mem[16'hEC19] = 8'h05;
mem[16'hEC1A] = 8'h9E;
mem[16'hEC1B] = 8'h85;
mem[16'hEC1C] = 8'h9E;
mem[16'hEC1D] = 8'h20;
mem[16'hEC1E] = 8'h07;
mem[16'hEC1F] = 8'hE9;
mem[16'hEC20] = 8'h84;
mem[16'hEC21] = 8'hA4;
mem[16'hEC22] = 8'h60;
mem[16'hEC23] = 8'hA5;
mem[16'hEC24] = 8'h9D;
mem[16'hEC25] = 8'hC9;
mem[16'hEC26] = 8'hA0;
mem[16'hEC27] = 8'hB0;
mem[16'hEC28] = 8'h20;
mem[16'hEC29] = 8'h20;
mem[16'hEC2A] = 8'hF2;
mem[16'hEC2B] = 8'hEB;
mem[16'hEC2C] = 8'h84;
mem[16'hEC2D] = 8'hAC;
mem[16'hEC2E] = 8'hA5;
mem[16'hEC2F] = 8'hA2;
mem[16'hEC30] = 8'h84;
mem[16'hEC31] = 8'hA2;
mem[16'hEC32] = 8'h49;
mem[16'hEC33] = 8'h80;
mem[16'hEC34] = 8'h2A;
mem[16'hEC35] = 8'hA9;
mem[16'hEC36] = 8'hA0;
mem[16'hEC37] = 8'h85;
mem[16'hEC38] = 8'h9D;
mem[16'hEC39] = 8'hA5;
mem[16'hEC3A] = 8'hA1;
mem[16'hEC3B] = 8'h85;
mem[16'hEC3C] = 8'h0D;
mem[16'hEC3D] = 8'h4C;
mem[16'hEC3E] = 8'h29;
mem[16'hEC3F] = 8'hE8;
mem[16'hEC40] = 8'h85;
mem[16'hEC41] = 8'h9E;
mem[16'hEC42] = 8'h85;
mem[16'hEC43] = 8'h9F;
mem[16'hEC44] = 8'h85;
mem[16'hEC45] = 8'hA0;
mem[16'hEC46] = 8'h85;
mem[16'hEC47] = 8'hA1;
mem[16'hEC48] = 8'hA8;
mem[16'hEC49] = 8'h60;
mem[16'hEC4A] = 8'hA0;
mem[16'hEC4B] = 8'h00;
mem[16'hEC4C] = 8'hA2;
mem[16'hEC4D] = 8'h0A;
mem[16'hEC4E] = 8'h94;
mem[16'hEC4F] = 8'h99;
mem[16'hEC50] = 8'hCA;
mem[16'hEC51] = 8'h10;
mem[16'hEC52] = 8'hFB;
mem[16'hEC53] = 8'h90;
mem[16'hEC54] = 8'h0F;
mem[16'hEC55] = 8'hC9;
mem[16'hEC56] = 8'h2D;
mem[16'hEC57] = 8'hD0;
mem[16'hEC58] = 8'h04;
mem[16'hEC59] = 8'h86;
mem[16'hEC5A] = 8'hA3;
mem[16'hEC5B] = 8'hF0;
mem[16'hEC5C] = 8'h04;
mem[16'hEC5D] = 8'hC9;
mem[16'hEC5E] = 8'h2B;
mem[16'hEC5F] = 8'hD0;
mem[16'hEC60] = 8'h05;
mem[16'hEC61] = 8'h20;
mem[16'hEC62] = 8'hB1;
mem[16'hEC63] = 8'h00;
mem[16'hEC64] = 8'h90;
mem[16'hEC65] = 8'h5B;
mem[16'hEC66] = 8'hC9;
mem[16'hEC67] = 8'h2E;
mem[16'hEC68] = 8'hF0;
mem[16'hEC69] = 8'h2E;
mem[16'hEC6A] = 8'hC9;
mem[16'hEC6B] = 8'h45;
mem[16'hEC6C] = 8'hD0;
mem[16'hEC6D] = 8'h30;
mem[16'hEC6E] = 8'h20;
mem[16'hEC6F] = 8'hB1;
mem[16'hEC70] = 8'h00;
mem[16'hEC71] = 8'h90;
mem[16'hEC72] = 8'h17;
mem[16'hEC73] = 8'hC9;
mem[16'hEC74] = 8'hC9;
mem[16'hEC75] = 8'hF0;
mem[16'hEC76] = 8'h0E;
mem[16'hEC77] = 8'hC9;
mem[16'hEC78] = 8'h2D;
mem[16'hEC79] = 8'hF0;
mem[16'hEC7A] = 8'h0A;
mem[16'hEC7B] = 8'hC9;
mem[16'hEC7C] = 8'hC8;
mem[16'hEC7D] = 8'hF0;
mem[16'hEC7E] = 8'h08;
mem[16'hEC7F] = 8'hC9;
mem[16'hEC80] = 8'h2B;
mem[16'hEC81] = 8'hF0;
mem[16'hEC82] = 8'h04;
mem[16'hEC83] = 8'hD0;
mem[16'hEC84] = 8'h07;
mem[16'hEC85] = 8'h66;
mem[16'hEC86] = 8'h9C;
mem[16'hEC87] = 8'h20;
mem[16'hEC88] = 8'hB1;
mem[16'hEC89] = 8'h00;
mem[16'hEC8A] = 8'h90;
mem[16'hEC8B] = 8'h5C;
mem[16'hEC8C] = 8'h24;
mem[16'hEC8D] = 8'h9C;
mem[16'hEC8E] = 8'h10;
mem[16'hEC8F] = 8'h0E;
mem[16'hEC90] = 8'hA9;
mem[16'hEC91] = 8'h00;
mem[16'hEC92] = 8'h38;
mem[16'hEC93] = 8'hE5;
mem[16'hEC94] = 8'h9A;
mem[16'hEC95] = 8'h4C;
mem[16'hEC96] = 8'hA0;
mem[16'hEC97] = 8'hEC;
mem[16'hEC98] = 8'h66;
mem[16'hEC99] = 8'h9B;
mem[16'hEC9A] = 8'h24;
mem[16'hEC9B] = 8'h9B;
mem[16'hEC9C] = 8'h50;
mem[16'hEC9D] = 8'hC3;
mem[16'hEC9E] = 8'hA5;
mem[16'hEC9F] = 8'h9A;
mem[16'hECA0] = 8'h38;
mem[16'hECA1] = 8'hE5;
mem[16'hECA2] = 8'h99;
mem[16'hECA3] = 8'h85;
mem[16'hECA4] = 8'h9A;
mem[16'hECA5] = 8'hF0;
mem[16'hECA6] = 8'h12;
mem[16'hECA7] = 8'h10;
mem[16'hECA8] = 8'h09;
mem[16'hECA9] = 8'h20;
mem[16'hECAA] = 8'h55;
mem[16'hECAB] = 8'hEA;
mem[16'hECAC] = 8'hE6;
mem[16'hECAD] = 8'h9A;
mem[16'hECAE] = 8'hD0;
mem[16'hECAF] = 8'hF9;
mem[16'hECB0] = 8'hF0;
mem[16'hECB1] = 8'h07;
mem[16'hECB2] = 8'h20;
mem[16'hECB3] = 8'h39;
mem[16'hECB4] = 8'hEA;
mem[16'hECB5] = 8'hC6;
mem[16'hECB6] = 8'h9A;
mem[16'hECB7] = 8'hD0;
mem[16'hECB8] = 8'hF9;
mem[16'hECB9] = 8'hA5;
mem[16'hECBA] = 8'hA3;
mem[16'hECBB] = 8'h30;
mem[16'hECBC] = 8'h01;
mem[16'hECBD] = 8'h60;
mem[16'hECBE] = 8'h4C;
mem[16'hECBF] = 8'hD0;
mem[16'hECC0] = 8'hEE;
mem[16'hECC1] = 8'h48;
mem[16'hECC2] = 8'h24;
mem[16'hECC3] = 8'h9B;
mem[16'hECC4] = 8'h10;
mem[16'hECC5] = 8'h02;
mem[16'hECC6] = 8'hE6;
mem[16'hECC7] = 8'h99;
mem[16'hECC8] = 8'h20;
mem[16'hECC9] = 8'h39;
mem[16'hECCA] = 8'hEA;
mem[16'hECCB] = 8'h68;
mem[16'hECCC] = 8'h38;
mem[16'hECCD] = 8'hE9;
mem[16'hECCE] = 8'h30;
mem[16'hECCF] = 8'h20;
mem[16'hECD0] = 8'hD5;
mem[16'hECD1] = 8'hEC;
mem[16'hECD2] = 8'h4C;
mem[16'hECD3] = 8'h61;
mem[16'hECD4] = 8'hEC;
mem[16'hECD5] = 8'h48;
mem[16'hECD6] = 8'h20;
mem[16'hECD7] = 8'h63;
mem[16'hECD8] = 8'hEB;
mem[16'hECD9] = 8'h68;
mem[16'hECDA] = 8'h20;
mem[16'hECDB] = 8'h93;
mem[16'hECDC] = 8'hEB;
mem[16'hECDD] = 8'hA5;
mem[16'hECDE] = 8'hAA;
mem[16'hECDF] = 8'h45;
mem[16'hECE0] = 8'hA2;
mem[16'hECE1] = 8'h85;
mem[16'hECE2] = 8'hAB;
mem[16'hECE3] = 8'hA6;
mem[16'hECE4] = 8'h9D;
mem[16'hECE5] = 8'h4C;
mem[16'hECE6] = 8'hC1;
mem[16'hECE7] = 8'hE7;
mem[16'hECE8] = 8'hA5;
mem[16'hECE9] = 8'h9A;
mem[16'hECEA] = 8'hC9;
mem[16'hECEB] = 8'h0A;
mem[16'hECEC] = 8'h90;
mem[16'hECED] = 8'h09;
mem[16'hECEE] = 8'hA9;
mem[16'hECEF] = 8'h64;
mem[16'hECF0] = 8'h24;
mem[16'hECF1] = 8'h9C;
mem[16'hECF2] = 8'h30;
mem[16'hECF3] = 8'h11;
mem[16'hECF4] = 8'h4C;
mem[16'hECF5] = 8'hD5;
mem[16'hECF6] = 8'hE8;
mem[16'hECF7] = 8'h0A;
mem[16'hECF8] = 8'h0A;
mem[16'hECF9] = 8'h18;
mem[16'hECFA] = 8'h65;
mem[16'hECFB] = 8'h9A;
mem[16'hECFC] = 8'h0A;
mem[16'hECFD] = 8'h18;
mem[16'hECFE] = 8'hA0;
mem[16'hECFF] = 8'h00;
mem[16'hED00] = 8'h71;
mem[16'hED01] = 8'hB8;
mem[16'hED02] = 8'h38;
mem[16'hED03] = 8'hE9;
mem[16'hED04] = 8'h30;
mem[16'hED05] = 8'h85;
mem[16'hED06] = 8'h9A;
mem[16'hED07] = 8'h4C;
mem[16'hED08] = 8'h87;
mem[16'hED09] = 8'hEC;
mem[16'hED0A] = 8'h9B;
mem[16'hED0B] = 8'h3E;
mem[16'hED0C] = 8'hBC;
mem[16'hED0D] = 8'h1F;
mem[16'hED0E] = 8'hFD;
mem[16'hED0F] = 8'h9E;
mem[16'hED10] = 8'h6E;
mem[16'hED11] = 8'h6B;
mem[16'hED12] = 8'h27;
mem[16'hED13] = 8'hFD;
mem[16'hED14] = 8'h9E;
mem[16'hED15] = 8'h6E;
mem[16'hED16] = 8'h6B;
mem[16'hED17] = 8'h28;
mem[16'hED18] = 8'h00;
mem[16'hED19] = 8'hA9;
mem[16'hED1A] = 8'h58;
mem[16'hED1B] = 8'hA0;
mem[16'hED1C] = 8'hD3;
mem[16'hED1D] = 8'h20;
mem[16'hED1E] = 8'h31;
mem[16'hED1F] = 8'hED;
mem[16'hED20] = 8'hA5;
mem[16'hED21] = 8'h76;
mem[16'hED22] = 8'hA6;
mem[16'hED23] = 8'h75;
mem[16'hED24] = 8'h85;
mem[16'hED25] = 8'h9E;
mem[16'hED26] = 8'h86;
mem[16'hED27] = 8'h9F;
mem[16'hED28] = 8'hA2;
mem[16'hED29] = 8'h90;
mem[16'hED2A] = 8'h38;
mem[16'hED2B] = 8'h20;
mem[16'hED2C] = 8'hA0;
mem[16'hED2D] = 8'hEB;
mem[16'hED2E] = 8'h20;
mem[16'hED2F] = 8'h34;
mem[16'hED30] = 8'hED;
mem[16'hED31] = 8'h4C;
mem[16'hED32] = 8'h3A;
mem[16'hED33] = 8'hDB;
mem[16'hED34] = 8'hA0;
mem[16'hED35] = 8'h01;
mem[16'hED36] = 8'hA9;
mem[16'hED37] = 8'h2D;
mem[16'hED38] = 8'h88;
mem[16'hED39] = 8'h24;
mem[16'hED3A] = 8'hA2;
mem[16'hED3B] = 8'h10;
mem[16'hED3C] = 8'h04;
mem[16'hED3D] = 8'hC8;
mem[16'hED3E] = 8'h99;
mem[16'hED3F] = 8'hFF;
mem[16'hED40] = 8'h00;
mem[16'hED41] = 8'h85;
mem[16'hED42] = 8'hA2;
mem[16'hED43] = 8'h84;
mem[16'hED44] = 8'hAD;
mem[16'hED45] = 8'hC8;
mem[16'hED46] = 8'hA9;
mem[16'hED47] = 8'h30;
mem[16'hED48] = 8'hA6;
mem[16'hED49] = 8'h9D;
mem[16'hED4A] = 8'hD0;
mem[16'hED4B] = 8'h03;
mem[16'hED4C] = 8'h4C;
mem[16'hED4D] = 8'h57;
mem[16'hED4E] = 8'hEE;
mem[16'hED4F] = 8'hA9;
mem[16'hED50] = 8'h00;
mem[16'hED51] = 8'hE0;
mem[16'hED52] = 8'h80;
mem[16'hED53] = 8'hF0;
mem[16'hED54] = 8'h02;
mem[16'hED55] = 8'hB0;
mem[16'hED56] = 8'h09;
mem[16'hED57] = 8'hA9;
mem[16'hED58] = 8'h14;
mem[16'hED59] = 8'hA0;
mem[16'hED5A] = 8'hED;
mem[16'hED5B] = 8'h20;
mem[16'hED5C] = 8'h7F;
mem[16'hED5D] = 8'hE9;
mem[16'hED5E] = 8'hA9;
mem[16'hED5F] = 8'hF7;
mem[16'hED60] = 8'h85;
mem[16'hED61] = 8'h99;
mem[16'hED62] = 8'hA9;
mem[16'hED63] = 8'h0F;
mem[16'hED64] = 8'hA0;
mem[16'hED65] = 8'hED;
mem[16'hED66] = 8'h20;
mem[16'hED67] = 8'hB2;
mem[16'hED68] = 8'hEB;
mem[16'hED69] = 8'hF0;
mem[16'hED6A] = 8'h1E;
mem[16'hED6B] = 8'h10;
mem[16'hED6C] = 8'h12;
mem[16'hED6D] = 8'hA9;
mem[16'hED6E] = 8'h0A;
mem[16'hED6F] = 8'hA0;
mem[16'hED70] = 8'hED;
mem[16'hED71] = 8'h20;
mem[16'hED72] = 8'hB2;
mem[16'hED73] = 8'hEB;
mem[16'hED74] = 8'hF0;
mem[16'hED75] = 8'h02;
mem[16'hED76] = 8'h10;
mem[16'hED77] = 8'h0E;
mem[16'hED78] = 8'h20;
mem[16'hED79] = 8'h39;
mem[16'hED7A] = 8'hEA;
mem[16'hED7B] = 8'hC6;
mem[16'hED7C] = 8'h99;
mem[16'hED7D] = 8'hD0;
mem[16'hED7E] = 8'hEE;
mem[16'hED7F] = 8'h20;
mem[16'hED80] = 8'h55;
mem[16'hED81] = 8'hEA;
mem[16'hED82] = 8'hE6;
mem[16'hED83] = 8'h99;
mem[16'hED84] = 8'hD0;
mem[16'hED85] = 8'hDC;
mem[16'hED86] = 8'h20;
mem[16'hED87] = 8'hA0;
mem[16'hED88] = 8'hE7;
mem[16'hED89] = 8'h20;
mem[16'hED8A] = 8'hF2;
mem[16'hED8B] = 8'hEB;
mem[16'hED8C] = 8'hA2;
mem[16'hED8D] = 8'h01;
mem[16'hED8E] = 8'hA5;
mem[16'hED8F] = 8'h99;
mem[16'hED90] = 8'h18;
mem[16'hED91] = 8'h69;
mem[16'hED92] = 8'h0A;
mem[16'hED93] = 8'h30;
mem[16'hED94] = 8'h09;
mem[16'hED95] = 8'hC9;
mem[16'hED96] = 8'h0B;
mem[16'hED97] = 8'hB0;
mem[16'hED98] = 8'h06;
mem[16'hED99] = 8'h69;
mem[16'hED9A] = 8'hFF;
mem[16'hED9B] = 8'hAA;
mem[16'hED9C] = 8'hA9;
mem[16'hED9D] = 8'h02;
mem[16'hED9E] = 8'h38;
mem[16'hED9F] = 8'hE9;
mem[16'hEDA0] = 8'h02;
mem[16'hEDA1] = 8'h85;
mem[16'hEDA2] = 8'h9A;
mem[16'hEDA3] = 8'h86;
mem[16'hEDA4] = 8'h99;
mem[16'hEDA5] = 8'h8A;
mem[16'hEDA6] = 8'hF0;
mem[16'hEDA7] = 8'h02;
mem[16'hEDA8] = 8'h10;
mem[16'hEDA9] = 8'h13;
mem[16'hEDAA] = 8'hA4;
mem[16'hEDAB] = 8'hAD;
mem[16'hEDAC] = 8'hA9;
mem[16'hEDAD] = 8'h2E;
mem[16'hEDAE] = 8'hC8;
mem[16'hEDAF] = 8'h99;
mem[16'hEDB0] = 8'hFF;
mem[16'hEDB1] = 8'h00;
mem[16'hEDB2] = 8'h8A;
mem[16'hEDB3] = 8'hF0;
mem[16'hEDB4] = 8'h06;
mem[16'hEDB5] = 8'hA9;
mem[16'hEDB6] = 8'h30;
mem[16'hEDB7] = 8'hC8;
mem[16'hEDB8] = 8'h99;
mem[16'hEDB9] = 8'hFF;
mem[16'hEDBA] = 8'h00;
mem[16'hEDBB] = 8'h84;
mem[16'hEDBC] = 8'hAD;
mem[16'hEDBD] = 8'hA0;
mem[16'hEDBE] = 8'h00;
mem[16'hEDBF] = 8'hA2;
mem[16'hEDC0] = 8'h80;
mem[16'hEDC1] = 8'hA5;
mem[16'hEDC2] = 8'hA1;
mem[16'hEDC3] = 8'h18;
mem[16'hEDC4] = 8'h79;
mem[16'hEDC5] = 8'h6C;
mem[16'hEDC6] = 8'hEE;
mem[16'hEDC7] = 8'h85;
mem[16'hEDC8] = 8'hA1;
mem[16'hEDC9] = 8'hA5;
mem[16'hEDCA] = 8'hA0;
mem[16'hEDCB] = 8'h79;
mem[16'hEDCC] = 8'h6B;
mem[16'hEDCD] = 8'hEE;
mem[16'hEDCE] = 8'h85;
mem[16'hEDCF] = 8'hA0;
mem[16'hEDD0] = 8'hA5;
mem[16'hEDD1] = 8'h9F;
mem[16'hEDD2] = 8'h79;
mem[16'hEDD3] = 8'h6A;
mem[16'hEDD4] = 8'hEE;
mem[16'hEDD5] = 8'h85;
mem[16'hEDD6] = 8'h9F;
mem[16'hEDD7] = 8'hA5;
mem[16'hEDD8] = 8'h9E;
mem[16'hEDD9] = 8'h79;
mem[16'hEDDA] = 8'h69;
mem[16'hEDDB] = 8'hEE;
mem[16'hEDDC] = 8'h85;
mem[16'hEDDD] = 8'h9E;
mem[16'hEDDE] = 8'hE8;
mem[16'hEDDF] = 8'hB0;
mem[16'hEDE0] = 8'h04;
mem[16'hEDE1] = 8'h10;
mem[16'hEDE2] = 8'hDE;
mem[16'hEDE3] = 8'h30;
mem[16'hEDE4] = 8'h02;
mem[16'hEDE5] = 8'h30;
mem[16'hEDE6] = 8'hDA;
mem[16'hEDE7] = 8'h8A;
mem[16'hEDE8] = 8'h90;
mem[16'hEDE9] = 8'h04;
mem[16'hEDEA] = 8'h49;
mem[16'hEDEB] = 8'hFF;
mem[16'hEDEC] = 8'h69;
mem[16'hEDED] = 8'h0A;
mem[16'hEDEE] = 8'h69;
mem[16'hEDEF] = 8'h2F;
mem[16'hEDF0] = 8'hC8;
mem[16'hEDF1] = 8'hC8;
mem[16'hEDF2] = 8'hC8;
mem[16'hEDF3] = 8'hC8;
mem[16'hEDF4] = 8'h84;
mem[16'hEDF5] = 8'h83;
mem[16'hEDF6] = 8'hA4;
mem[16'hEDF7] = 8'hAD;
mem[16'hEDF8] = 8'hC8;
mem[16'hEDF9] = 8'hAA;
mem[16'hEDFA] = 8'h29;
mem[16'hEDFB] = 8'h7F;
mem[16'hEDFC] = 8'h99;
mem[16'hEDFD] = 8'hFF;
mem[16'hEDFE] = 8'h00;
mem[16'hEDFF] = 8'hC6;
mem[16'hEE00] = 8'h99;
mem[16'hEE01] = 8'hD0;
mem[16'hEE02] = 8'h06;
mem[16'hEE03] = 8'hA9;
mem[16'hEE04] = 8'h2E;
mem[16'hEE05] = 8'hC8;
mem[16'hEE06] = 8'h99;
mem[16'hEE07] = 8'hFF;
mem[16'hEE08] = 8'h00;
mem[16'hEE09] = 8'h84;
mem[16'hEE0A] = 8'hAD;
mem[16'hEE0B] = 8'hA4;
mem[16'hEE0C] = 8'h83;
mem[16'hEE0D] = 8'h8A;
mem[16'hEE0E] = 8'h49;
mem[16'hEE0F] = 8'hFF;
mem[16'hEE10] = 8'h29;
mem[16'hEE11] = 8'h80;
mem[16'hEE12] = 8'hAA;
mem[16'hEE13] = 8'hC0;
mem[16'hEE14] = 8'h24;
mem[16'hEE15] = 8'hD0;
mem[16'hEE16] = 8'hAA;
mem[16'hEE17] = 8'hA4;
mem[16'hEE18] = 8'hAD;
mem[16'hEE19] = 8'hB9;
mem[16'hEE1A] = 8'hFF;
mem[16'hEE1B] = 8'h00;
mem[16'hEE1C] = 8'h88;
mem[16'hEE1D] = 8'hC9;
mem[16'hEE1E] = 8'h30;
mem[16'hEE1F] = 8'hF0;
mem[16'hEE20] = 8'hF8;
mem[16'hEE21] = 8'hC9;
mem[16'hEE22] = 8'h2E;
mem[16'hEE23] = 8'hF0;
mem[16'hEE24] = 8'h01;
mem[16'hEE25] = 8'hC8;
mem[16'hEE26] = 8'hA9;
mem[16'hEE27] = 8'h2B;
mem[16'hEE28] = 8'hA6;
mem[16'hEE29] = 8'h9A;
mem[16'hEE2A] = 8'hF0;
mem[16'hEE2B] = 8'h2E;
mem[16'hEE2C] = 8'h10;
mem[16'hEE2D] = 8'h08;
mem[16'hEE2E] = 8'hA9;
mem[16'hEE2F] = 8'h00;
mem[16'hEE30] = 8'h38;
mem[16'hEE31] = 8'hE5;
mem[16'hEE32] = 8'h9A;
mem[16'hEE33] = 8'hAA;
mem[16'hEE34] = 8'hA9;
mem[16'hEE35] = 8'h2D;
mem[16'hEE36] = 8'h99;
mem[16'hEE37] = 8'h01;
mem[16'hEE38] = 8'h01;
mem[16'hEE39] = 8'hA9;
mem[16'hEE3A] = 8'h45;
mem[16'hEE3B] = 8'h99;
mem[16'hEE3C] = 8'h00;
mem[16'hEE3D] = 8'h01;
mem[16'hEE3E] = 8'h8A;
mem[16'hEE3F] = 8'hA2;
mem[16'hEE40] = 8'h2F;
mem[16'hEE41] = 8'h38;
mem[16'hEE42] = 8'hE8;
mem[16'hEE43] = 8'hE9;
mem[16'hEE44] = 8'h0A;
mem[16'hEE45] = 8'hB0;
mem[16'hEE46] = 8'hFB;
mem[16'hEE47] = 8'h69;
mem[16'hEE48] = 8'h3A;
mem[16'hEE49] = 8'h99;
mem[16'hEE4A] = 8'h03;
mem[16'hEE4B] = 8'h01;
mem[16'hEE4C] = 8'h8A;
mem[16'hEE4D] = 8'h99;
mem[16'hEE4E] = 8'h02;
mem[16'hEE4F] = 8'h01;
mem[16'hEE50] = 8'hA9;
mem[16'hEE51] = 8'h00;
mem[16'hEE52] = 8'h99;
mem[16'hEE53] = 8'h04;
mem[16'hEE54] = 8'h01;
mem[16'hEE55] = 8'hF0;
mem[16'hEE56] = 8'h08;
mem[16'hEE57] = 8'h99;
mem[16'hEE58] = 8'hFF;
mem[16'hEE59] = 8'h00;
mem[16'hEE5A] = 8'hA9;
mem[16'hEE5B] = 8'h00;
mem[16'hEE5C] = 8'h99;
mem[16'hEE5D] = 8'h00;
mem[16'hEE5E] = 8'h01;
mem[16'hEE5F] = 8'hA9;
mem[16'hEE60] = 8'h00;
mem[16'hEE61] = 8'hA0;
mem[16'hEE62] = 8'h01;
mem[16'hEE63] = 8'h60;
mem[16'hEE64] = 8'h80;
mem[16'hEE65] = 8'h00;
mem[16'hEE66] = 8'h00;
mem[16'hEE67] = 8'h00;
mem[16'hEE68] = 8'h00;
mem[16'hEE69] = 8'hFA;
mem[16'hEE6A] = 8'h0A;
mem[16'hEE6B] = 8'h1F;
mem[16'hEE6C] = 8'h00;
mem[16'hEE6D] = 8'h00;
mem[16'hEE6E] = 8'h98;
mem[16'hEE6F] = 8'h96;
mem[16'hEE70] = 8'h80;
mem[16'hEE71] = 8'hFF;
mem[16'hEE72] = 8'hF0;
mem[16'hEE73] = 8'hBD;
mem[16'hEE74] = 8'hC0;
mem[16'hEE75] = 8'h00;
mem[16'hEE76] = 8'h01;
mem[16'hEE77] = 8'h86;
mem[16'hEE78] = 8'hA0;
mem[16'hEE79] = 8'hFF;
mem[16'hEE7A] = 8'hFF;
mem[16'hEE7B] = 8'hD8;
mem[16'hEE7C] = 8'hF0;
mem[16'hEE7D] = 8'h00;
mem[16'hEE7E] = 8'h00;
mem[16'hEE7F] = 8'h03;
mem[16'hEE80] = 8'hE8;
mem[16'hEE81] = 8'hFF;
mem[16'hEE82] = 8'hFF;
mem[16'hEE83] = 8'hFF;
mem[16'hEE84] = 8'h9C;
mem[16'hEE85] = 8'h00;
mem[16'hEE86] = 8'h00;
mem[16'hEE87] = 8'h00;
mem[16'hEE88] = 8'h0A;
mem[16'hEE89] = 8'hFF;
mem[16'hEE8A] = 8'hFF;
mem[16'hEE8B] = 8'hFF;
mem[16'hEE8C] = 8'hFF;
mem[16'hEE8D] = 8'h20;
mem[16'hEE8E] = 8'h63;
mem[16'hEE8F] = 8'hEB;
mem[16'hEE90] = 8'hA9;
mem[16'hEE91] = 8'h64;
mem[16'hEE92] = 8'hA0;
mem[16'hEE93] = 8'hEE;
mem[16'hEE94] = 8'h20;
mem[16'hEE95] = 8'hF9;
mem[16'hEE96] = 8'hEA;
mem[16'hEE97] = 8'hF0;
mem[16'hEE98] = 8'h70;
mem[16'hEE99] = 8'hA5;
mem[16'hEE9A] = 8'hA5;
mem[16'hEE9B] = 8'hD0;
mem[16'hEE9C] = 8'h03;
mem[16'hEE9D] = 8'h4C;
mem[16'hEE9E] = 8'h50;
mem[16'hEE9F] = 8'hE8;
mem[16'hEEA0] = 8'hA2;
mem[16'hEEA1] = 8'h8A;
mem[16'hEEA2] = 8'hA0;
mem[16'hEEA3] = 8'h00;
mem[16'hEEA4] = 8'h20;
mem[16'hEEA5] = 8'h2B;
mem[16'hEEA6] = 8'hEB;
mem[16'hEEA7] = 8'hA5;
mem[16'hEEA8] = 8'hAA;
mem[16'hEEA9] = 8'h10;
mem[16'hEEAA] = 8'h0F;
mem[16'hEEAB] = 8'h20;
mem[16'hEEAC] = 8'h23;
mem[16'hEEAD] = 8'hEC;
mem[16'hEEAE] = 8'hA9;
mem[16'hEEAF] = 8'h8A;
mem[16'hEEB0] = 8'hA0;
mem[16'hEEB1] = 8'h00;
mem[16'hEEB2] = 8'h20;
mem[16'hEEB3] = 8'hB2;
mem[16'hEEB4] = 8'hEB;
mem[16'hEEB5] = 8'hD0;
mem[16'hEEB6] = 8'h03;
mem[16'hEEB7] = 8'h98;
mem[16'hEEB8] = 8'hA4;
mem[16'hEEB9] = 8'h0D;
mem[16'hEEBA] = 8'h20;
mem[16'hEEBB] = 8'h55;
mem[16'hEEBC] = 8'hEB;
mem[16'hEEBD] = 8'h98;
mem[16'hEEBE] = 8'h48;
mem[16'hEEBF] = 8'h20;
mem[16'hEEC0] = 8'h41;
mem[16'hEEC1] = 8'hE9;
mem[16'hEEC2] = 8'hA9;
mem[16'hEEC3] = 8'h8A;
mem[16'hEEC4] = 8'hA0;
mem[16'hEEC5] = 8'h00;
mem[16'hEEC6] = 8'h20;
mem[16'hEEC7] = 8'h7F;
mem[16'hEEC8] = 8'hE9;
mem[16'hEEC9] = 8'h20;
mem[16'hEECA] = 8'h09;
mem[16'hEECB] = 8'hEF;
mem[16'hEECC] = 8'h68;
mem[16'hEECD] = 8'h4A;
mem[16'hEECE] = 8'h90;
mem[16'hEECF] = 8'h0A;
mem[16'hEED0] = 8'hA5;
mem[16'hEED1] = 8'h9D;
mem[16'hEED2] = 8'hF0;
mem[16'hEED3] = 8'h06;
mem[16'hEED4] = 8'hA5;
mem[16'hEED5] = 8'hA2;
mem[16'hEED6] = 8'h49;
mem[16'hEED7] = 8'hFF;
mem[16'hEED8] = 8'h85;
mem[16'hEED9] = 8'hA2;
mem[16'hEEDA] = 8'h60;
mem[16'hEEDB] = 8'h81;
mem[16'hEEDC] = 8'h38;
mem[16'hEEDD] = 8'hAA;
mem[16'hEEDE] = 8'h3B;
mem[16'hEEDF] = 8'h29;
mem[16'hEEE0] = 8'h07;
mem[16'hEEE1] = 8'h71;
mem[16'hEEE2] = 8'h34;
mem[16'hEEE3] = 8'h58;
mem[16'hEEE4] = 8'h3E;
mem[16'hEEE5] = 8'h56;
mem[16'hEEE6] = 8'h74;
mem[16'hEEE7] = 8'h16;
mem[16'hEEE8] = 8'h7E;
mem[16'hEEE9] = 8'hB3;
mem[16'hEEEA] = 8'h1B;
mem[16'hEEEB] = 8'h77;
mem[16'hEEEC] = 8'h2F;
mem[16'hEEED] = 8'hEE;
mem[16'hEEEE] = 8'hE3;
mem[16'hEEEF] = 8'h85;
mem[16'hEEF0] = 8'h7A;
mem[16'hEEF1] = 8'h1D;
mem[16'hEEF2] = 8'h84;
mem[16'hEEF3] = 8'h1C;
mem[16'hEEF4] = 8'h2A;
mem[16'hEEF5] = 8'h7C;
mem[16'hEEF6] = 8'h63;
mem[16'hEEF7] = 8'h59;
mem[16'hEEF8] = 8'h58;
mem[16'hEEF9] = 8'h0A;
mem[16'hEEFA] = 8'h7E;
mem[16'hEEFB] = 8'h75;
mem[16'hEEFC] = 8'hFD;
mem[16'hEEFD] = 8'hE7;
mem[16'hEEFE] = 8'hC6;
mem[16'hEEFF] = 8'h80;
mem[16'hEF00] = 8'h31;
mem[16'hEF01] = 8'h72;
mem[16'hEF02] = 8'h18;
mem[16'hEF03] = 8'h10;
mem[16'hEF04] = 8'h81;
mem[16'hEF05] = 8'h00;
mem[16'hEF06] = 8'h00;
mem[16'hEF07] = 8'h00;
mem[16'hEF08] = 8'h00;
mem[16'hEF09] = 8'hA9;
mem[16'hEF0A] = 8'hDB;
mem[16'hEF0B] = 8'hA0;
mem[16'hEF0C] = 8'hEE;
mem[16'hEF0D] = 8'h20;
mem[16'hEF0E] = 8'h7F;
mem[16'hEF0F] = 8'hE9;
mem[16'hEF10] = 8'hA5;
mem[16'hEF11] = 8'hAC;
mem[16'hEF12] = 8'h69;
mem[16'hEF13] = 8'h50;
mem[16'hEF14] = 8'h90;
mem[16'hEF15] = 8'h03;
mem[16'hEF16] = 8'h20;
mem[16'hEF17] = 8'h7A;
mem[16'hEF18] = 8'hEB;
mem[16'hEF19] = 8'h85;
mem[16'hEF1A] = 8'h92;
mem[16'hEF1B] = 8'h20;
mem[16'hEF1C] = 8'h66;
mem[16'hEF1D] = 8'hEB;
mem[16'hEF1E] = 8'hA5;
mem[16'hEF1F] = 8'h9D;
mem[16'hEF20] = 8'hC9;
mem[16'hEF21] = 8'h88;
mem[16'hEF22] = 8'h90;
mem[16'hEF23] = 8'h03;
mem[16'hEF24] = 8'h20;
mem[16'hEF25] = 8'h2B;
mem[16'hEF26] = 8'hEA;
mem[16'hEF27] = 8'h20;
mem[16'hEF28] = 8'h23;
mem[16'hEF29] = 8'hEC;
mem[16'hEF2A] = 8'hA5;
mem[16'hEF2B] = 8'h0D;
mem[16'hEF2C] = 8'h18;
mem[16'hEF2D] = 8'h69;
mem[16'hEF2E] = 8'h81;
mem[16'hEF2F] = 8'hF0;
mem[16'hEF30] = 8'hF3;
mem[16'hEF31] = 8'h38;
mem[16'hEF32] = 8'hE9;
mem[16'hEF33] = 8'h01;
mem[16'hEF34] = 8'h48;
mem[16'hEF35] = 8'hA2;
mem[16'hEF36] = 8'h05;
mem[16'hEF37] = 8'hB5;
mem[16'hEF38] = 8'hA5;
mem[16'hEF39] = 8'hB4;
mem[16'hEF3A] = 8'h9D;
mem[16'hEF3B] = 8'h95;
mem[16'hEF3C] = 8'h9D;
mem[16'hEF3D] = 8'h94;
mem[16'hEF3E] = 8'hA5;
mem[16'hEF3F] = 8'hCA;
mem[16'hEF40] = 8'h10;
mem[16'hEF41] = 8'hF5;
mem[16'hEF42] = 8'hA5;
mem[16'hEF43] = 8'h92;
mem[16'hEF44] = 8'h85;
mem[16'hEF45] = 8'hAC;
mem[16'hEF46] = 8'h20;
mem[16'hEF47] = 8'hAA;
mem[16'hEF48] = 8'hE7;
mem[16'hEF49] = 8'h20;
mem[16'hEF4A] = 8'hD0;
mem[16'hEF4B] = 8'hEE;
mem[16'hEF4C] = 8'hA9;
mem[16'hEF4D] = 8'hE0;
mem[16'hEF4E] = 8'hA0;
mem[16'hEF4F] = 8'hEE;
mem[16'hEF50] = 8'h20;
mem[16'hEF51] = 8'h72;
mem[16'hEF52] = 8'hEF;
mem[16'hEF53] = 8'hA9;
mem[16'hEF54] = 8'h00;
mem[16'hEF55] = 8'h85;
mem[16'hEF56] = 8'hAB;
mem[16'hEF57] = 8'h68;
mem[16'hEF58] = 8'h20;
mem[16'hEF59] = 8'h10;
mem[16'hEF5A] = 8'hEA;
mem[16'hEF5B] = 8'h60;
mem[16'hEF5C] = 8'h85;
mem[16'hEF5D] = 8'hAD;
mem[16'hEF5E] = 8'h84;
mem[16'hEF5F] = 8'hAE;
mem[16'hEF60] = 8'h20;
mem[16'hEF61] = 8'h21;
mem[16'hEF62] = 8'hEB;
mem[16'hEF63] = 8'hA9;
mem[16'hEF64] = 8'h93;
mem[16'hEF65] = 8'h20;
mem[16'hEF66] = 8'h7F;
mem[16'hEF67] = 8'hE9;
mem[16'hEF68] = 8'h20;
mem[16'hEF69] = 8'h76;
mem[16'hEF6A] = 8'hEF;
mem[16'hEF6B] = 8'hA9;
mem[16'hEF6C] = 8'h93;
mem[16'hEF6D] = 8'hA0;
mem[16'hEF6E] = 8'h00;
mem[16'hEF6F] = 8'h4C;
mem[16'hEF70] = 8'h7F;
mem[16'hEF71] = 8'hE9;
mem[16'hEF72] = 8'h85;
mem[16'hEF73] = 8'hAD;
mem[16'hEF74] = 8'h84;
mem[16'hEF75] = 8'hAE;
mem[16'hEF76] = 8'h20;
mem[16'hEF77] = 8'h1E;
mem[16'hEF78] = 8'hEB;
mem[16'hEF79] = 8'hB1;
mem[16'hEF7A] = 8'hAD;
mem[16'hEF7B] = 8'h85;
mem[16'hEF7C] = 8'hA3;
mem[16'hEF7D] = 8'hA4;
mem[16'hEF7E] = 8'hAD;
mem[16'hEF7F] = 8'hC8;
mem[16'hEF80] = 8'h98;
mem[16'hEF81] = 8'hD0;
mem[16'hEF82] = 8'h02;
mem[16'hEF83] = 8'hE6;
mem[16'hEF84] = 8'hAE;
mem[16'hEF85] = 8'h85;
mem[16'hEF86] = 8'hAD;
mem[16'hEF87] = 8'hA4;
mem[16'hEF88] = 8'hAE;
mem[16'hEF89] = 8'h20;
mem[16'hEF8A] = 8'h7F;
mem[16'hEF8B] = 8'hE9;
mem[16'hEF8C] = 8'hA5;
mem[16'hEF8D] = 8'hAD;
mem[16'hEF8E] = 8'hA4;
mem[16'hEF8F] = 8'hAE;
mem[16'hEF90] = 8'h18;
mem[16'hEF91] = 8'h69;
mem[16'hEF92] = 8'h05;
mem[16'hEF93] = 8'h90;
mem[16'hEF94] = 8'h01;
mem[16'hEF95] = 8'hC8;
mem[16'hEF96] = 8'h85;
mem[16'hEF97] = 8'hAD;
mem[16'hEF98] = 8'h84;
mem[16'hEF99] = 8'hAE;
mem[16'hEF9A] = 8'h20;
mem[16'hEF9B] = 8'hBE;
mem[16'hEF9C] = 8'hE7;
mem[16'hEF9D] = 8'hA9;
mem[16'hEF9E] = 8'h98;
mem[16'hEF9F] = 8'hA0;
mem[16'hEFA0] = 8'h00;
mem[16'hEFA1] = 8'hC6;
mem[16'hEFA2] = 8'hA3;
mem[16'hEFA3] = 8'hD0;
mem[16'hEFA4] = 8'hE4;
mem[16'hEFA5] = 8'h60;
mem[16'hEFA6] = 8'h98;
mem[16'hEFA7] = 8'h35;
mem[16'hEFA8] = 8'h44;
mem[16'hEFA9] = 8'h7A;
mem[16'hEFAA] = 8'h68;
mem[16'hEFAB] = 8'h28;
mem[16'hEFAC] = 8'hB1;
mem[16'hEFAD] = 8'h46;
mem[16'hEFAE] = 8'h20;
mem[16'hEFAF] = 8'h82;
mem[16'hEFB0] = 8'hEB;
mem[16'hEFB1] = 8'hAA;
mem[16'hEFB2] = 8'h30;
mem[16'hEFB3] = 8'h18;
mem[16'hEFB4] = 8'hA9;
mem[16'hEFB5] = 8'hC9;
mem[16'hEFB6] = 8'hA0;
mem[16'hEFB7] = 8'h00;
mem[16'hEFB8] = 8'h20;
mem[16'hEFB9] = 8'hF9;
mem[16'hEFBA] = 8'hEA;
mem[16'hEFBB] = 8'h8A;
mem[16'hEFBC] = 8'hF0;
mem[16'hEFBD] = 8'hE7;
mem[16'hEFBE] = 8'hA9;
mem[16'hEFBF] = 8'hA6;
mem[16'hEFC0] = 8'hA0;
mem[16'hEFC1] = 8'hEF;
mem[16'hEFC2] = 8'h20;
mem[16'hEFC3] = 8'h7F;
mem[16'hEFC4] = 8'hE9;
mem[16'hEFC5] = 8'hA9;
mem[16'hEFC6] = 8'hAA;
mem[16'hEFC7] = 8'hA0;
mem[16'hEFC8] = 8'hEF;
mem[16'hEFC9] = 8'h20;
mem[16'hEFCA] = 8'hBE;
mem[16'hEFCB] = 8'hE7;
mem[16'hEFCC] = 8'hA6;
mem[16'hEFCD] = 8'hA1;
mem[16'hEFCE] = 8'hA5;
mem[16'hEFCF] = 8'h9E;
mem[16'hEFD0] = 8'h85;
mem[16'hEFD1] = 8'hA1;
mem[16'hEFD2] = 8'h86;
mem[16'hEFD3] = 8'h9E;
mem[16'hEFD4] = 8'hA9;
mem[16'hEFD5] = 8'h00;
mem[16'hEFD6] = 8'h85;
mem[16'hEFD7] = 8'hA2;
mem[16'hEFD8] = 8'hA5;
mem[16'hEFD9] = 8'h9D;
mem[16'hEFDA] = 8'h85;
mem[16'hEFDB] = 8'hAC;
mem[16'hEFDC] = 8'hA9;
mem[16'hEFDD] = 8'h80;
mem[16'hEFDE] = 8'h85;
mem[16'hEFDF] = 8'h9D;
mem[16'hEFE0] = 8'h20;
mem[16'hEFE1] = 8'h2E;
mem[16'hEFE2] = 8'hE8;
mem[16'hEFE3] = 8'hA2;
mem[16'hEFE4] = 8'hC9;
mem[16'hEFE5] = 8'hA0;
mem[16'hEFE6] = 8'h00;
mem[16'hEFE7] = 8'h4C;
mem[16'hEFE8] = 8'h2B;
mem[16'hEFE9] = 8'hEB;
mem[16'hEFEA] = 8'hA9;
mem[16'hEFEB] = 8'h66;
mem[16'hEFEC] = 8'hA0;
mem[16'hEFED] = 8'hF0;
mem[16'hEFEE] = 8'h20;
mem[16'hEFEF] = 8'hBE;
mem[16'hEFF0] = 8'hE7;
mem[16'hEFF1] = 8'h20;
mem[16'hEFF2] = 8'h63;
mem[16'hEFF3] = 8'hEB;
mem[16'hEFF4] = 8'hA9;
mem[16'hEFF5] = 8'h6B;
mem[16'hEFF6] = 8'hA0;
mem[16'hEFF7] = 8'hF0;
mem[16'hEFF8] = 8'hA6;
mem[16'hEFF9] = 8'hAA;
mem[16'hEFFA] = 8'h20;
mem[16'hEFFB] = 8'h5E;
mem[16'hEFFC] = 8'hEA;
mem[16'hEFFD] = 8'h20;
mem[16'hEFFE] = 8'h63;
mem[16'hEFFF] = 8'hEB;
mem[16'hF000] = 8'h20;
mem[16'hF001] = 8'h23;
mem[16'hF002] = 8'hEC;
mem[16'hF003] = 8'hA9;
mem[16'hF004] = 8'h00;
mem[16'hF005] = 8'h85;
mem[16'hF006] = 8'hAB;
mem[16'hF007] = 8'h20;
mem[16'hF008] = 8'hAA;
mem[16'hF009] = 8'hE7;
mem[16'hF00A] = 8'hA9;
mem[16'hF00B] = 8'h70;
mem[16'hF00C] = 8'hA0;
mem[16'hF00D] = 8'hF0;
mem[16'hF00E] = 8'h20;
mem[16'hF00F] = 8'hA7;
mem[16'hF010] = 8'hE7;
mem[16'hF011] = 8'hA5;
mem[16'hF012] = 8'hA2;
mem[16'hF013] = 8'h48;
mem[16'hF014] = 8'h10;
mem[16'hF015] = 8'h0D;
mem[16'hF016] = 8'h20;
mem[16'hF017] = 8'hA0;
mem[16'hF018] = 8'hE7;
mem[16'hF019] = 8'hA5;
mem[16'hF01A] = 8'hA2;
mem[16'hF01B] = 8'h30;
mem[16'hF01C] = 8'h09;
mem[16'hF01D] = 8'hA5;
mem[16'hF01E] = 8'h16;
mem[16'hF01F] = 8'h49;
mem[16'hF020] = 8'hFF;
mem[16'hF021] = 8'h85;
mem[16'hF022] = 8'h16;
mem[16'hF023] = 8'h20;
mem[16'hF024] = 8'hD0;
mem[16'hF025] = 8'hEE;
mem[16'hF026] = 8'hA9;
mem[16'hF027] = 8'h70;
mem[16'hF028] = 8'hA0;
mem[16'hF029] = 8'hF0;
mem[16'hF02A] = 8'h20;
mem[16'hF02B] = 8'hBE;
mem[16'hF02C] = 8'hE7;
mem[16'hF02D] = 8'h68;
mem[16'hF02E] = 8'h10;
mem[16'hF02F] = 8'h03;
mem[16'hF030] = 8'h20;
mem[16'hF031] = 8'hD0;
mem[16'hF032] = 8'hEE;
mem[16'hF033] = 8'hA9;
mem[16'hF034] = 8'h75;
mem[16'hF035] = 8'hA0;
mem[16'hF036] = 8'hF0;
mem[16'hF037] = 8'h4C;
mem[16'hF038] = 8'h5C;
mem[16'hF039] = 8'hEF;
mem[16'hF03A] = 8'h20;
mem[16'hF03B] = 8'h21;
mem[16'hF03C] = 8'hEB;
mem[16'hF03D] = 8'hA9;
mem[16'hF03E] = 8'h00;
mem[16'hF03F] = 8'h85;
mem[16'hF040] = 8'h16;
mem[16'hF041] = 8'h20;
mem[16'hF042] = 8'hF1;
mem[16'hF043] = 8'hEF;
mem[16'hF044] = 8'hA2;
mem[16'hF045] = 8'h8A;
mem[16'hF046] = 8'hA0;
mem[16'hF047] = 8'h00;
mem[16'hF048] = 8'h20;
mem[16'hF049] = 8'hE7;
mem[16'hF04A] = 8'hEF;
mem[16'hF04B] = 8'hA9;
mem[16'hF04C] = 8'h93;
mem[16'hF04D] = 8'hA0;
mem[16'hF04E] = 8'h00;
mem[16'hF04F] = 8'h20;
mem[16'hF050] = 8'hF9;
mem[16'hF051] = 8'hEA;
mem[16'hF052] = 8'hA9;
mem[16'hF053] = 8'h00;
mem[16'hF054] = 8'h85;
mem[16'hF055] = 8'hA2;
mem[16'hF056] = 8'hA5;
mem[16'hF057] = 8'h16;
mem[16'hF058] = 8'h20;
mem[16'hF059] = 8'h62;
mem[16'hF05A] = 8'hF0;
mem[16'hF05B] = 8'hA9;
mem[16'hF05C] = 8'h8A;
mem[16'hF05D] = 8'hA0;
mem[16'hF05E] = 8'h00;
mem[16'hF05F] = 8'h4C;
mem[16'hF060] = 8'h66;
mem[16'hF061] = 8'hEA;
mem[16'hF062] = 8'h48;
mem[16'hF063] = 8'h4C;
mem[16'hF064] = 8'h23;
mem[16'hF065] = 8'hF0;
mem[16'hF066] = 8'h81;
mem[16'hF067] = 8'h49;
mem[16'hF068] = 8'h0F;
mem[16'hF069] = 8'hDA;
mem[16'hF06A] = 8'hA2;
mem[16'hF06B] = 8'h83;
mem[16'hF06C] = 8'h49;
mem[16'hF06D] = 8'h0F;
mem[16'hF06E] = 8'hDA;
mem[16'hF06F] = 8'hA2;
mem[16'hF070] = 8'h7F;
mem[16'hF071] = 8'h00;
mem[16'hF072] = 8'h00;
mem[16'hF073] = 8'h00;
mem[16'hF074] = 8'h00;
mem[16'hF075] = 8'h05;
mem[16'hF076] = 8'h84;
mem[16'hF077] = 8'hE6;
mem[16'hF078] = 8'h1A;
mem[16'hF079] = 8'h2D;
mem[16'hF07A] = 8'h1B;
mem[16'hF07B] = 8'h86;
mem[16'hF07C] = 8'h28;
mem[16'hF07D] = 8'h07;
mem[16'hF07E] = 8'hFB;
mem[16'hF07F] = 8'hF8;
mem[16'hF080] = 8'h87;
mem[16'hF081] = 8'h99;
mem[16'hF082] = 8'h68;
mem[16'hF083] = 8'h89;
mem[16'hF084] = 8'h01;
mem[16'hF085] = 8'h87;
mem[16'hF086] = 8'h23;
mem[16'hF087] = 8'h35;
mem[16'hF088] = 8'hDF;
mem[16'hF089] = 8'hE1;
mem[16'hF08A] = 8'h86;
mem[16'hF08B] = 8'hA5;
mem[16'hF08C] = 8'h5D;
mem[16'hF08D] = 8'hE7;
mem[16'hF08E] = 8'h28;
mem[16'hF08F] = 8'h83;
mem[16'hF090] = 8'h49;
mem[16'hF091] = 8'h0F;
mem[16'hF092] = 8'hDA;
mem[16'hF093] = 8'hA2;
mem[16'hF094] = 8'hA6;
mem[16'hF095] = 8'hD3;
mem[16'hF096] = 8'hC1;
mem[16'hF097] = 8'hC8;
mem[16'hF098] = 8'hD4;
mem[16'hF099] = 8'hC8;
mem[16'hF09A] = 8'hD5;
mem[16'hF09B] = 8'hC4;
mem[16'hF09C] = 8'hCE;
mem[16'hF09D] = 8'hCA;
mem[16'hF09E] = 8'hA5;
mem[16'hF09F] = 8'hA2;
mem[16'hF0A0] = 8'h48;
mem[16'hF0A1] = 8'h10;
mem[16'hF0A2] = 8'h03;
mem[16'hF0A3] = 8'h20;
mem[16'hF0A4] = 8'hD0;
mem[16'hF0A5] = 8'hEE;
mem[16'hF0A6] = 8'hA5;
mem[16'hF0A7] = 8'h9D;
mem[16'hF0A8] = 8'h48;
mem[16'hF0A9] = 8'hC9;
mem[16'hF0AA] = 8'h81;
mem[16'hF0AB] = 8'h90;
mem[16'hF0AC] = 8'h07;
mem[16'hF0AD] = 8'hA9;
mem[16'hF0AE] = 8'h13;
mem[16'hF0AF] = 8'hA0;
mem[16'hF0B0] = 8'hE9;
mem[16'hF0B1] = 8'h20;
mem[16'hF0B2] = 8'h66;
mem[16'hF0B3] = 8'hEA;
mem[16'hF0B4] = 8'hA9;
mem[16'hF0B5] = 8'hCE;
mem[16'hF0B6] = 8'hA0;
mem[16'hF0B7] = 8'hF0;
mem[16'hF0B8] = 8'h20;
mem[16'hF0B9] = 8'h5C;
mem[16'hF0BA] = 8'hEF;
mem[16'hF0BB] = 8'h68;
mem[16'hF0BC] = 8'hC9;
mem[16'hF0BD] = 8'h81;
mem[16'hF0BE] = 8'h90;
mem[16'hF0BF] = 8'h07;
mem[16'hF0C0] = 8'hA9;
mem[16'hF0C1] = 8'h66;
mem[16'hF0C2] = 8'hA0;
mem[16'hF0C3] = 8'hF0;
mem[16'hF0C4] = 8'h20;
mem[16'hF0C5] = 8'hA7;
mem[16'hF0C6] = 8'hE7;
mem[16'hF0C7] = 8'h68;
mem[16'hF0C8] = 8'h10;
mem[16'hF0C9] = 8'h03;
mem[16'hF0CA] = 8'h4C;
mem[16'hF0CB] = 8'hD0;
mem[16'hF0CC] = 8'hEE;
mem[16'hF0CD] = 8'h60;
mem[16'hF0CE] = 8'h0B;
mem[16'hF0CF] = 8'h76;
mem[16'hF0D0] = 8'hB3;
mem[16'hF0D1] = 8'h83;
mem[16'hF0D2] = 8'hBD;
mem[16'hF0D3] = 8'hD3;
mem[16'hF0D4] = 8'h79;
mem[16'hF0D5] = 8'h1E;
mem[16'hF0D6] = 8'hF4;
mem[16'hF0D7] = 8'hA6;
mem[16'hF0D8] = 8'hF5;
mem[16'hF0D9] = 8'h7B;
mem[16'hF0DA] = 8'h83;
mem[16'hF0DB] = 8'hFC;
mem[16'hF0DC] = 8'hB0;
mem[16'hF0DD] = 8'h10;
mem[16'hF0DE] = 8'h7C;
mem[16'hF0DF] = 8'h0C;
mem[16'hF0E0] = 8'h1F;
mem[16'hF0E1] = 8'h67;
mem[16'hF0E2] = 8'hCA;
mem[16'hF0E3] = 8'h7C;
mem[16'hF0E4] = 8'hDE;
mem[16'hF0E5] = 8'h53;
mem[16'hF0E6] = 8'hCB;
mem[16'hF0E7] = 8'hC1;
mem[16'hF0E8] = 8'h7D;
mem[16'hF0E9] = 8'h14;
mem[16'hF0EA] = 8'h64;
mem[16'hF0EB] = 8'h70;
mem[16'hF0EC] = 8'h4C;
mem[16'hF0ED] = 8'h7D;
mem[16'hF0EE] = 8'hB7;
mem[16'hF0EF] = 8'hEA;
mem[16'hF0F0] = 8'h51;
mem[16'hF0F1] = 8'h7A;
mem[16'hF0F2] = 8'h7D;
mem[16'hF0F3] = 8'h63;
mem[16'hF0F4] = 8'h30;
mem[16'hF0F5] = 8'h88;
mem[16'hF0F6] = 8'h7E;
mem[16'hF0F7] = 8'h7E;
mem[16'hF0F8] = 8'h92;
mem[16'hF0F9] = 8'h44;
mem[16'hF0FA] = 8'h99;
mem[16'hF0FB] = 8'h3A;
mem[16'hF0FC] = 8'h7E;
mem[16'hF0FD] = 8'h4C;
mem[16'hF0FE] = 8'hCC;
mem[16'hF0FF] = 8'h91;
mem[16'hF100] = 8'hC7;
mem[16'hF101] = 8'h7F;
mem[16'hF102] = 8'hAA;
mem[16'hF103] = 8'hAA;
mem[16'hF104] = 8'hAA;
mem[16'hF105] = 8'h13;
mem[16'hF106] = 8'h81;
mem[16'hF107] = 8'h00;
mem[16'hF108] = 8'h00;
mem[16'hF109] = 8'h00;
mem[16'hF10A] = 8'h00;
mem[16'hF10B] = 8'hE6;
mem[16'hF10C] = 8'hB8;
mem[16'hF10D] = 8'hD0;
mem[16'hF10E] = 8'h02;
mem[16'hF10F] = 8'hE6;
mem[16'hF110] = 8'hB9;
mem[16'hF111] = 8'hAD;
mem[16'hF112] = 8'h60;
mem[16'hF113] = 8'hEA;
mem[16'hF114] = 8'hC9;
mem[16'hF115] = 8'h3A;
mem[16'hF116] = 8'hB0;
mem[16'hF117] = 8'h0A;
mem[16'hF118] = 8'hC9;
mem[16'hF119] = 8'h20;
mem[16'hF11A] = 8'hF0;
mem[16'hF11B] = 8'hEF;
mem[16'hF11C] = 8'h38;
mem[16'hF11D] = 8'hE9;
mem[16'hF11E] = 8'h30;
mem[16'hF11F] = 8'h38;
mem[16'hF120] = 8'hE9;
mem[16'hF121] = 8'hD0;
mem[16'hF122] = 8'h60;
mem[16'hF123] = 8'h80;
mem[16'hF124] = 8'h4F;
mem[16'hF125] = 8'hC7;
mem[16'hF126] = 8'h52;
mem[16'hF127] = 8'h58;
mem[16'hF128] = 8'hA2;
mem[16'hF129] = 8'hFF;
mem[16'hF12A] = 8'h86;
mem[16'hF12B] = 8'h76;
mem[16'hF12C] = 8'hA2;
mem[16'hF12D] = 8'hFB;
mem[16'hF12E] = 8'h9A;
mem[16'hF12F] = 8'hA9;
mem[16'hF130] = 8'h28;
mem[16'hF131] = 8'hA0;
mem[16'hF132] = 8'hF1;
mem[16'hF133] = 8'h85;
mem[16'hF134] = 8'h01;
mem[16'hF135] = 8'h84;
mem[16'hF136] = 8'h02;
mem[16'hF137] = 8'h85;
mem[16'hF138] = 8'h04;
mem[16'hF139] = 8'h84;
mem[16'hF13A] = 8'h05;
mem[16'hF13B] = 8'h20;
mem[16'hF13C] = 8'h73;
mem[16'hF13D] = 8'hF2;
mem[16'hF13E] = 8'hA9;
mem[16'hF13F] = 8'h4C;
mem[16'hF140] = 8'h85;
mem[16'hF141] = 8'h00;
mem[16'hF142] = 8'h85;
mem[16'hF143] = 8'h03;
mem[16'hF144] = 8'h85;
mem[16'hF145] = 8'h90;
mem[16'hF146] = 8'h85;
mem[16'hF147] = 8'h0A;
mem[16'hF148] = 8'hA9;
mem[16'hF149] = 8'h99;
mem[16'hF14A] = 8'hA0;
mem[16'hF14B] = 8'hE1;
mem[16'hF14C] = 8'h85;
mem[16'hF14D] = 8'h0B;
mem[16'hF14E] = 8'h84;
mem[16'hF14F] = 8'h0C;
mem[16'hF150] = 8'hA2;
mem[16'hF151] = 8'h1C;
mem[16'hF152] = 8'hBD;
mem[16'hF153] = 8'h0A;
mem[16'hF154] = 8'hF1;
mem[16'hF155] = 8'h95;
mem[16'hF156] = 8'hB0;
mem[16'hF157] = 8'h86;
mem[16'hF158] = 8'hF1;
mem[16'hF159] = 8'hCA;
mem[16'hF15A] = 8'hD0;
mem[16'hF15B] = 8'hF6;
mem[16'hF15C] = 8'h86;
mem[16'hF15D] = 8'hF2;
mem[16'hF15E] = 8'h8A;
mem[16'hF15F] = 8'h85;
mem[16'hF160] = 8'hA4;
mem[16'hF161] = 8'h85;
mem[16'hF162] = 8'h54;
mem[16'hF163] = 8'h48;
mem[16'hF164] = 8'hA9;
mem[16'hF165] = 8'h03;
mem[16'hF166] = 8'h85;
mem[16'hF167] = 8'h8F;
mem[16'hF168] = 8'h20;
mem[16'hF169] = 8'hFB;
mem[16'hF16A] = 8'hDA;
mem[16'hF16B] = 8'hA9;
mem[16'hF16C] = 8'h01;
mem[16'hF16D] = 8'h8D;
mem[16'hF16E] = 8'hFD;
mem[16'hF16F] = 8'h01;
mem[16'hF170] = 8'h8D;
mem[16'hF171] = 8'hFC;
mem[16'hF172] = 8'h01;
mem[16'hF173] = 8'hA2;
mem[16'hF174] = 8'h55;
mem[16'hF175] = 8'h86;
mem[16'hF176] = 8'h52;
mem[16'hF177] = 8'hA9;
mem[16'hF178] = 8'h00;
mem[16'hF179] = 8'hA0;
mem[16'hF17A] = 8'h08;
mem[16'hF17B] = 8'h85;
mem[16'hF17C] = 8'h50;
mem[16'hF17D] = 8'h84;
mem[16'hF17E] = 8'h51;
mem[16'hF17F] = 8'hA0;
mem[16'hF180] = 8'h00;
mem[16'hF181] = 8'hE6;
mem[16'hF182] = 8'h51;
mem[16'hF183] = 8'hB1;
mem[16'hF184] = 8'h50;
mem[16'hF185] = 8'h49;
mem[16'hF186] = 8'hFF;
mem[16'hF187] = 8'h91;
mem[16'hF188] = 8'h50;
mem[16'hF189] = 8'hD1;
mem[16'hF18A] = 8'h50;
mem[16'hF18B] = 8'hD0;
mem[16'hF18C] = 8'h08;
mem[16'hF18D] = 8'h49;
mem[16'hF18E] = 8'hFF;
mem[16'hF18F] = 8'h91;
mem[16'hF190] = 8'h50;
mem[16'hF191] = 8'hD1;
mem[16'hF192] = 8'h50;
mem[16'hF193] = 8'hF0;
mem[16'hF194] = 8'hEC;
mem[16'hF195] = 8'hA4;
mem[16'hF196] = 8'h50;
mem[16'hF197] = 8'hA5;
mem[16'hF198] = 8'h51;
mem[16'hF199] = 8'h29;
mem[16'hF19A] = 8'hF0;
mem[16'hF19B] = 8'h84;
mem[16'hF19C] = 8'h73;
mem[16'hF19D] = 8'h85;
mem[16'hF19E] = 8'h74;
mem[16'hF19F] = 8'h84;
mem[16'hF1A0] = 8'h6F;
mem[16'hF1A1] = 8'h85;
mem[16'hF1A2] = 8'h70;
mem[16'hF1A3] = 8'hA2;
mem[16'hF1A4] = 8'h00;
mem[16'hF1A5] = 8'hA0;
mem[16'hF1A6] = 8'h08;
mem[16'hF1A7] = 8'h86;
mem[16'hF1A8] = 8'h67;
mem[16'hF1A9] = 8'h84;
mem[16'hF1AA] = 8'h68;
mem[16'hF1AB] = 8'hA0;
mem[16'hF1AC] = 8'h00;
mem[16'hF1AD] = 8'h84;
mem[16'hF1AE] = 8'hD6;
mem[16'hF1AF] = 8'h98;
mem[16'hF1B0] = 8'h91;
mem[16'hF1B1] = 8'h67;
mem[16'hF1B2] = 8'hE6;
mem[16'hF1B3] = 8'h67;
mem[16'hF1B4] = 8'hD0;
mem[16'hF1B5] = 8'h02;
mem[16'hF1B6] = 8'hE6;
mem[16'hF1B7] = 8'h68;
mem[16'hF1B8] = 8'hA5;
mem[16'hF1B9] = 8'h67;
mem[16'hF1BA] = 8'hA4;
mem[16'hF1BB] = 8'h68;
mem[16'hF1BC] = 8'h20;
mem[16'hF1BD] = 8'hE3;
mem[16'hF1BE] = 8'hD3;
mem[16'hF1BF] = 8'h20;
mem[16'hF1C0] = 8'h4B;
mem[16'hF1C1] = 8'hD6;
mem[16'hF1C2] = 8'hA9;
mem[16'hF1C3] = 8'h3A;
mem[16'hF1C4] = 8'hA0;
mem[16'hF1C5] = 8'hDB;
mem[16'hF1C6] = 8'h85;
mem[16'hF1C7] = 8'h04;
mem[16'hF1C8] = 8'h84;
mem[16'hF1C9] = 8'h05;
mem[16'hF1CA] = 8'hA9;
mem[16'hF1CB] = 8'h3C;
mem[16'hF1CC] = 8'hA0;
mem[16'hF1CD] = 8'hD4;
mem[16'hF1CE] = 8'h85;
mem[16'hF1CF] = 8'h01;
mem[16'hF1D0] = 8'h84;
mem[16'hF1D1] = 8'h02;
mem[16'hF1D2] = 8'h6C;
mem[16'hF1D3] = 8'h01;
mem[16'hF1D4] = 8'h00;
mem[16'hF1D5] = 8'h20;
mem[16'hF1D6] = 8'h67;
mem[16'hF1D7] = 8'hDD;
mem[16'hF1D8] = 8'h20;
mem[16'hF1D9] = 8'h52;
mem[16'hF1DA] = 8'hE7;
mem[16'hF1DB] = 8'h6C;
mem[16'hF1DC] = 8'h50;
mem[16'hF1DD] = 8'h00;
mem[16'hF1DE] = 8'h20;
mem[16'hF1DF] = 8'hF8;
mem[16'hF1E0] = 8'hE6;
mem[16'hF1E1] = 8'h8A;
mem[16'hF1E2] = 8'h4C;
mem[16'hF1E3] = 8'h8B;
mem[16'hF1E4] = 8'hFE;
mem[16'hF1E5] = 8'h20;
mem[16'hF1E6] = 8'hF8;
mem[16'hF1E7] = 8'hE6;
mem[16'hF1E8] = 8'h8A;
mem[16'hF1E9] = 8'h4C;
mem[16'hF1EA] = 8'h95;
mem[16'hF1EB] = 8'hFE;
mem[16'hF1EC] = 8'h20;
mem[16'hF1ED] = 8'hF8;
mem[16'hF1EE] = 8'hE6;
mem[16'hF1EF] = 8'hE0;
mem[16'hF1F0] = 8'h30;
mem[16'hF1F1] = 8'hB0;
mem[16'hF1F2] = 8'h13;
mem[16'hF1F3] = 8'h86;
mem[16'hF1F4] = 8'hF0;
mem[16'hF1F5] = 8'hA9;
mem[16'hF1F6] = 8'h2C;
mem[16'hF1F7] = 8'h20;
mem[16'hF1F8] = 8'hC0;
mem[16'hF1F9] = 8'hDE;
mem[16'hF1FA] = 8'h20;
mem[16'hF1FB] = 8'hF8;
mem[16'hF1FC] = 8'hE6;
mem[16'hF1FD] = 8'hE0;
mem[16'hF1FE] = 8'h30;
mem[16'hF1FF] = 8'hB0;
mem[16'hF200] = 8'h05;
mem[16'hF201] = 8'h86;
mem[16'hF202] = 8'h2C;
mem[16'hF203] = 8'h86;
mem[16'hF204] = 8'h2D;
mem[16'hF205] = 8'h60;
mem[16'hF206] = 8'h4C;
mem[16'hF207] = 8'h99;
mem[16'hF208] = 8'hE1;
mem[16'hF209] = 8'h20;
mem[16'hF20A] = 8'hEC;
mem[16'hF20B] = 8'hF1;
mem[16'hF20C] = 8'hE4;
mem[16'hF20D] = 8'hF0;
mem[16'hF20E] = 8'hB0;
mem[16'hF20F] = 8'h08;
mem[16'hF210] = 8'hA5;
mem[16'hF211] = 8'hF0;
mem[16'hF212] = 8'h85;
mem[16'hF213] = 8'h2C;
mem[16'hF214] = 8'h85;
mem[16'hF215] = 8'h2D;
mem[16'hF216] = 8'h86;
mem[16'hF217] = 8'hF0;
mem[16'hF218] = 8'hA9;
mem[16'hF219] = 8'hC5;
mem[16'hF21A] = 8'h20;
mem[16'hF21B] = 8'hC0;
mem[16'hF21C] = 8'hDE;
mem[16'hF21D] = 8'h20;
mem[16'hF21E] = 8'hF8;
mem[16'hF21F] = 8'hE6;
mem[16'hF220] = 8'hE0;
mem[16'hF221] = 8'h30;
mem[16'hF222] = 8'hB0;
mem[16'hF223] = 8'hE2;
mem[16'hF224] = 8'h60;
mem[16'hF225] = 8'h20;
mem[16'hF226] = 8'hEC;
mem[16'hF227] = 8'hF1;
mem[16'hF228] = 8'h8A;
mem[16'hF229] = 8'hA4;
mem[16'hF22A] = 8'hF0;
mem[16'hF22B] = 8'hC0;
mem[16'hF22C] = 8'h28;
mem[16'hF22D] = 8'hB0;
mem[16'hF22E] = 8'hD7;
mem[16'hF22F] = 8'h4C;
mem[16'hF230] = 8'h00;
mem[16'hF231] = 8'hF8;
mem[16'hF232] = 8'h20;
mem[16'hF233] = 8'h09;
mem[16'hF234] = 8'hF2;
mem[16'hF235] = 8'h8A;
mem[16'hF236] = 8'hA4;
mem[16'hF237] = 8'h2C;
mem[16'hF238] = 8'hC0;
mem[16'hF239] = 8'h28;
mem[16'hF23A] = 8'hB0;
mem[16'hF23B] = 8'hCA;
mem[16'hF23C] = 8'hA4;
mem[16'hF23D] = 8'hF0;
mem[16'hF23E] = 8'h4C;
mem[16'hF23F] = 8'h19;
mem[16'hF240] = 8'hF8;
mem[16'hF241] = 8'h20;
mem[16'hF242] = 8'h09;
mem[16'hF243] = 8'hF2;
mem[16'hF244] = 8'h8A;
mem[16'hF245] = 8'hA8;
mem[16'hF246] = 8'hC0;
mem[16'hF247] = 8'h28;
mem[16'hF248] = 8'hB0;
mem[16'hF249] = 8'hBC;
mem[16'hF24A] = 8'hA5;
mem[16'hF24B] = 8'hF0;
mem[16'hF24C] = 8'h4C;
mem[16'hF24D] = 8'h28;
mem[16'hF24E] = 8'hF8;
mem[16'hF24F] = 8'h20;
mem[16'hF250] = 8'hF8;
mem[16'hF251] = 8'hE6;
mem[16'hF252] = 8'h8A;
mem[16'hF253] = 8'h4C;
mem[16'hF254] = 8'h64;
mem[16'hF255] = 8'hF8;
mem[16'hF256] = 8'h20;
mem[16'hF257] = 8'hF8;
mem[16'hF258] = 8'hE6;
mem[16'hF259] = 8'hCA;
mem[16'hF25A] = 8'h8A;
mem[16'hF25B] = 8'hC9;
mem[16'hF25C] = 8'h18;
mem[16'hF25D] = 8'hB0;
mem[16'hF25E] = 8'hA7;
mem[16'hF25F] = 8'h4C;
mem[16'hF260] = 8'h5B;
mem[16'hF261] = 8'hFB;
mem[16'hF262] = 8'h20;
mem[16'hF263] = 8'hF8;
mem[16'hF264] = 8'hE6;
mem[16'hF265] = 8'h8A;
mem[16'hF266] = 8'h49;
mem[16'hF267] = 8'hFF;
mem[16'hF268] = 8'hAA;
mem[16'hF269] = 8'hE8;
mem[16'hF26A] = 8'h86;
mem[16'hF26B] = 8'hF1;
mem[16'hF26C] = 8'h60;
mem[16'hF26D] = 8'h38;
mem[16'hF26E] = 8'h90;
mem[16'hF26F] = 8'h18;
mem[16'hF270] = 8'h66;
mem[16'hF271] = 8'hF2;
mem[16'hF272] = 8'h60;
mem[16'hF273] = 8'hA9;
mem[16'hF274] = 8'hFF;
mem[16'hF275] = 8'hD0;
mem[16'hF276] = 8'h02;
mem[16'hF277] = 8'hA9;
mem[16'hF278] = 8'h3F;
mem[16'hF279] = 8'hA2;
mem[16'hF27A] = 8'h00;
mem[16'hF27B] = 8'h85;
mem[16'hF27C] = 8'h32;
mem[16'hF27D] = 8'h86;
mem[16'hF27E] = 8'hF3;
mem[16'hF27F] = 8'h60;
mem[16'hF280] = 8'hA9;
mem[16'hF281] = 8'h7F;
mem[16'hF282] = 8'hA2;
mem[16'hF283] = 8'h40;
mem[16'hF284] = 8'hD0;
mem[16'hF285] = 8'hF5;
mem[16'hF286] = 8'h20;
mem[16'hF287] = 8'h67;
mem[16'hF288] = 8'hDD;
mem[16'hF289] = 8'h20;
mem[16'hF28A] = 8'h52;
mem[16'hF28B] = 8'hE7;
mem[16'hF28C] = 8'hA5;
mem[16'hF28D] = 8'h50;
mem[16'hF28E] = 8'hC5;
mem[16'hF28F] = 8'h6D;
mem[16'hF290] = 8'hA5;
mem[16'hF291] = 8'h51;
mem[16'hF292] = 8'hE5;
mem[16'hF293] = 8'h6E;
mem[16'hF294] = 8'hB0;
mem[16'hF295] = 8'h03;
mem[16'hF296] = 8'h4C;
mem[16'hF297] = 8'h10;
mem[16'hF298] = 8'hD4;
mem[16'hF299] = 8'hA5;
mem[16'hF29A] = 8'h50;
mem[16'hF29B] = 8'h85;
mem[16'hF29C] = 8'h73;
mem[16'hF29D] = 8'h85;
mem[16'hF29E] = 8'h6F;
mem[16'hF29F] = 8'hA5;
mem[16'hF2A0] = 8'h51;
mem[16'hF2A1] = 8'h85;
mem[16'hF2A2] = 8'h74;
mem[16'hF2A3] = 8'h85;
mem[16'hF2A4] = 8'h70;
mem[16'hF2A5] = 8'h60;
mem[16'hF2A6] = 8'h20;
mem[16'hF2A7] = 8'h67;
mem[16'hF2A8] = 8'hDD;
mem[16'hF2A9] = 8'h20;
mem[16'hF2AA] = 8'h52;
mem[16'hF2AB] = 8'hE7;
mem[16'hF2AC] = 8'hA5;
mem[16'hF2AD] = 8'h50;
mem[16'hF2AE] = 8'hC5;
mem[16'hF2AF] = 8'h73;
mem[16'hF2B0] = 8'hA5;
mem[16'hF2B1] = 8'h51;
mem[16'hF2B2] = 8'hE5;
mem[16'hF2B3] = 8'h74;
mem[16'hF2B4] = 8'hB0;
mem[16'hF2B5] = 8'hE0;
mem[16'hF2B6] = 8'hA5;
mem[16'hF2B7] = 8'h50;
mem[16'hF2B8] = 8'hC5;
mem[16'hF2B9] = 8'h69;
mem[16'hF2BA] = 8'hA5;
mem[16'hF2BB] = 8'h51;
mem[16'hF2BC] = 8'hE5;
mem[16'hF2BD] = 8'h6A;
mem[16'hF2BE] = 8'h90;
mem[16'hF2BF] = 8'hD6;
mem[16'hF2C0] = 8'hA5;
mem[16'hF2C1] = 8'h50;
mem[16'hF2C2] = 8'h85;
mem[16'hF2C3] = 8'h69;
mem[16'hF2C4] = 8'hA5;
mem[16'hF2C5] = 8'h51;
mem[16'hF2C6] = 8'h85;
mem[16'hF2C7] = 8'h6A;
mem[16'hF2C8] = 8'h4C;
mem[16'hF2C9] = 8'h6C;
mem[16'hF2CA] = 8'hD6;
mem[16'hF2CB] = 8'hA9;
mem[16'hF2CC] = 8'hAB;
mem[16'hF2CD] = 8'h20;
mem[16'hF2CE] = 8'hC0;
mem[16'hF2CF] = 8'hDE;
mem[16'hF2D0] = 8'hA5;
mem[16'hF2D1] = 8'hB8;
mem[16'hF2D2] = 8'h85;
mem[16'hF2D3] = 8'hF4;
mem[16'hF2D4] = 8'hA5;
mem[16'hF2D5] = 8'hB9;
mem[16'hF2D6] = 8'h85;
mem[16'hF2D7] = 8'hF5;
mem[16'hF2D8] = 8'h38;
mem[16'hF2D9] = 8'h66;
mem[16'hF2DA] = 8'hD8;
mem[16'hF2DB] = 8'hA5;
mem[16'hF2DC] = 8'h75;
mem[16'hF2DD] = 8'h85;
mem[16'hF2DE] = 8'hF6;
mem[16'hF2DF] = 8'hA5;
mem[16'hF2E0] = 8'h76;
mem[16'hF2E1] = 8'h85;
mem[16'hF2E2] = 8'hF7;
mem[16'hF2E3] = 8'h20;
mem[16'hF2E4] = 8'hA6;
mem[16'hF2E5] = 8'hD9;
mem[16'hF2E6] = 8'h4C;
mem[16'hF2E7] = 8'h98;
mem[16'hF2E8] = 8'hD9;
mem[16'hF2E9] = 8'h86;
mem[16'hF2EA] = 8'hDE;
mem[16'hF2EB] = 8'hA6;
mem[16'hF2EC] = 8'hF8;
mem[16'hF2ED] = 8'h86;
mem[16'hF2EE] = 8'hDF;
mem[16'hF2EF] = 8'hA5;
mem[16'hF2F0] = 8'h75;
mem[16'hF2F1] = 8'h85;
mem[16'hF2F2] = 8'hDA;
mem[16'hF2F3] = 8'hA5;
mem[16'hF2F4] = 8'h76;
mem[16'hF2F5] = 8'h85;
mem[16'hF2F6] = 8'hDB;
mem[16'hF2F7] = 8'hA5;
mem[16'hF2F8] = 8'h79;
mem[16'hF2F9] = 8'h85;
mem[16'hF2FA] = 8'hDC;
mem[16'hF2FB] = 8'hA5;
mem[16'hF2FC] = 8'h7A;
mem[16'hF2FD] = 8'h85;
mem[16'hF2FE] = 8'hDD;
mem[16'hF2FF] = 8'hA5;
mem[16'hF300] = 8'hF4;
mem[16'hF301] = 8'h85;
mem[16'hF302] = 8'hB8;
mem[16'hF303] = 8'hA5;
mem[16'hF304] = 8'hF5;
mem[16'hF305] = 8'h85;
mem[16'hF306] = 8'hB9;
mem[16'hF307] = 8'hA5;
mem[16'hF308] = 8'hF6;
mem[16'hF309] = 8'h85;
mem[16'hF30A] = 8'h75;
mem[16'hF30B] = 8'hA5;
mem[16'hF30C] = 8'hF7;
mem[16'hF30D] = 8'h85;
mem[16'hF30E] = 8'h76;
mem[16'hF30F] = 8'h20;
mem[16'hF310] = 8'hB7;
mem[16'hF311] = 8'h00;
mem[16'hF312] = 8'h20;
mem[16'hF313] = 8'h3E;
mem[16'hF314] = 8'hD9;
mem[16'hF315] = 8'h4C;
mem[16'hF316] = 8'hD2;
mem[16'hF317] = 8'hD7;
mem[16'hF318] = 8'hA5;
mem[16'hF319] = 8'hDA;
mem[16'hF31A] = 8'h85;
mem[16'hF31B] = 8'h75;
mem[16'hF31C] = 8'hA5;
mem[16'hF31D] = 8'hDB;
mem[16'hF31E] = 8'h85;
mem[16'hF31F] = 8'h76;
mem[16'hF320] = 8'hA5;
mem[16'hF321] = 8'hDC;
mem[16'hF322] = 8'h85;
mem[16'hF323] = 8'hB8;
mem[16'hF324] = 8'hA5;
mem[16'hF325] = 8'hDD;
mem[16'hF326] = 8'h85;
mem[16'hF327] = 8'hB9;
mem[16'hF328] = 8'hA6;
mem[16'hF329] = 8'hDF;
mem[16'hF32A] = 8'h9A;
mem[16'hF32B] = 8'h4C;
mem[16'hF32C] = 8'hD2;
mem[16'hF32D] = 8'hD7;
mem[16'hF32E] = 8'h4C;
mem[16'hF32F] = 8'hC9;
mem[16'hF330] = 8'hDE;
mem[16'hF331] = 8'hB0;
mem[16'hF332] = 8'hFB;
mem[16'hF333] = 8'hA6;
mem[16'hF334] = 8'hAF;
mem[16'hF335] = 8'h86;
mem[16'hF336] = 8'h69;
mem[16'hF337] = 8'hA6;
mem[16'hF338] = 8'hB0;
mem[16'hF339] = 8'h86;
mem[16'hF33A] = 8'h6A;
mem[16'hF33B] = 8'h20;
mem[16'hF33C] = 8'h0C;
mem[16'hF33D] = 8'hDA;
mem[16'hF33E] = 8'h20;
mem[16'hF33F] = 8'h1A;
mem[16'hF340] = 8'hD6;
mem[16'hF341] = 8'hA5;
mem[16'hF342] = 8'h9B;
mem[16'hF343] = 8'h85;
mem[16'hF344] = 8'h60;
mem[16'hF345] = 8'hA5;
mem[16'hF346] = 8'h9C;
mem[16'hF347] = 8'h85;
mem[16'hF348] = 8'h61;
mem[16'hF349] = 8'hA9;
mem[16'hF34A] = 8'h2C;
mem[16'hF34B] = 8'h20;
mem[16'hF34C] = 8'hC0;
mem[16'hF34D] = 8'hDE;
mem[16'hF34E] = 8'h20;
mem[16'hF34F] = 8'h0C;
mem[16'hF350] = 8'hDA;
mem[16'hF351] = 8'hE6;
mem[16'hF352] = 8'h50;
mem[16'hF353] = 8'hD0;
mem[16'hF354] = 8'h02;
mem[16'hF355] = 8'hE6;
mem[16'hF356] = 8'h51;
mem[16'hF357] = 8'h20;
mem[16'hF358] = 8'h1A;
mem[16'hF359] = 8'hD6;
mem[16'hF35A] = 8'hA5;
mem[16'hF35B] = 8'h9B;
mem[16'hF35C] = 8'hC5;
mem[16'hF35D] = 8'h60;
mem[16'hF35E] = 8'hA5;
mem[16'hF35F] = 8'h9C;
mem[16'hF360] = 8'hE5;
mem[16'hF361] = 8'h61;
mem[16'hF362] = 8'hB0;
mem[16'hF363] = 8'h01;
mem[16'hF364] = 8'h60;
mem[16'hF365] = 8'hA0;
mem[16'hF366] = 8'h00;
mem[16'hF367] = 8'hB1;
mem[16'hF368] = 8'h9B;
mem[16'hF369] = 8'h91;
mem[16'hF36A] = 8'h60;
mem[16'hF36B] = 8'hE6;
mem[16'hF36C] = 8'h9B;
mem[16'hF36D] = 8'hD0;
mem[16'hF36E] = 8'h02;
mem[16'hF36F] = 8'hE6;
mem[16'hF370] = 8'h9C;
mem[16'hF371] = 8'hE6;
mem[16'hF372] = 8'h60;
mem[16'hF373] = 8'hD0;
mem[16'hF374] = 8'h02;
mem[16'hF375] = 8'hE6;
mem[16'hF376] = 8'h61;
mem[16'hF377] = 8'hA5;
mem[16'hF378] = 8'h69;
mem[16'hF379] = 8'hC5;
mem[16'hF37A] = 8'h9B;
mem[16'hF37B] = 8'hA5;
mem[16'hF37C] = 8'h6A;
mem[16'hF37D] = 8'hE5;
mem[16'hF37E] = 8'h9C;
mem[16'hF37F] = 8'hB0;
mem[16'hF380] = 8'hE6;
mem[16'hF381] = 8'hA6;
mem[16'hF382] = 8'h61;
mem[16'hF383] = 8'hA4;
mem[16'hF384] = 8'h60;
mem[16'hF385] = 8'hD0;
mem[16'hF386] = 8'h01;
mem[16'hF387] = 8'hCA;
mem[16'hF388] = 8'h88;
mem[16'hF389] = 8'h86;
mem[16'hF38A] = 8'h6A;
mem[16'hF38B] = 8'h84;
mem[16'hF38C] = 8'h69;
mem[16'hF38D] = 8'h4C;
mem[16'hF38E] = 8'hF2;
mem[16'hF38F] = 8'hD4;
mem[16'hF390] = 8'hAD;
mem[16'hF391] = 8'h56;
mem[16'hF392] = 8'hC0;
mem[16'hF393] = 8'hAD;
mem[16'hF394] = 8'h53;
mem[16'hF395] = 8'hC0;
mem[16'hF396] = 8'h4C;
mem[16'hF397] = 8'h40;
mem[16'hF398] = 8'hFB;
mem[16'hF399] = 8'hAD;
mem[16'hF39A] = 8'h54;
mem[16'hF39B] = 8'hC0;
mem[16'hF39C] = 8'h4C;
mem[16'hF39D] = 8'h39;
mem[16'hF39E] = 8'hFB;
mem[16'hF39F] = 8'h20;
mem[16'hF3A0] = 8'hD9;
mem[16'hF3A1] = 8'hF7;
mem[16'hF3A2] = 8'hA0;
mem[16'hF3A3] = 8'h03;
mem[16'hF3A4] = 8'hB1;
mem[16'hF3A5] = 8'h9B;
mem[16'hF3A6] = 8'hAA;
mem[16'hF3A7] = 8'h88;
mem[16'hF3A8] = 8'hB1;
mem[16'hF3A9] = 8'h9B;
mem[16'hF3AA] = 8'hE9;
mem[16'hF3AB] = 8'h01;
mem[16'hF3AC] = 8'hB0;
mem[16'hF3AD] = 8'h01;
mem[16'hF3AE] = 8'hCA;
mem[16'hF3AF] = 8'h85;
mem[16'hF3B0] = 8'h50;
mem[16'hF3B1] = 8'h86;
mem[16'hF3B2] = 8'h51;
mem[16'hF3B3] = 8'h20;
mem[16'hF3B4] = 8'hCD;
mem[16'hF3B5] = 8'hFE;
mem[16'hF3B6] = 8'h20;
mem[16'hF3B7] = 8'hBC;
mem[16'hF3B8] = 8'hF7;
mem[16'hF3B9] = 8'h4C;
mem[16'hF3BA] = 8'hCD;
mem[16'hF3BB] = 8'hFE;
mem[16'hF3BC] = 8'h20;
mem[16'hF3BD] = 8'hD9;
mem[16'hF3BE] = 8'hF7;
mem[16'hF3BF] = 8'h20;
mem[16'hF3C0] = 8'hFD;
mem[16'hF3C1] = 8'hFE;
mem[16'hF3C2] = 8'hA0;
mem[16'hF3C3] = 8'h02;
mem[16'hF3C4] = 8'hB1;
mem[16'hF3C5] = 8'h9B;
mem[16'hF3C6] = 8'hC5;
mem[16'hF3C7] = 8'h50;
mem[16'hF3C8] = 8'hC8;
mem[16'hF3C9] = 8'hB1;
mem[16'hF3CA] = 8'h9B;
mem[16'hF3CB] = 8'hE5;
mem[16'hF3CC] = 8'h51;
mem[16'hF3CD] = 8'hB0;
mem[16'hF3CE] = 8'h03;
mem[16'hF3CF] = 8'h4C;
mem[16'hF3D0] = 8'h10;
mem[16'hF3D1] = 8'hD4;
mem[16'hF3D2] = 8'h20;
mem[16'hF3D3] = 8'hBC;
mem[16'hF3D4] = 8'hF7;
mem[16'hF3D5] = 8'h4C;
mem[16'hF3D6] = 8'hFD;
mem[16'hF3D7] = 8'hFE;
mem[16'hF3D8] = 8'h2C;
mem[16'hF3D9] = 8'h55;
mem[16'hF3DA] = 8'hC0;
mem[16'hF3DB] = 8'h2C;
mem[16'hF3DC] = 8'h52;
mem[16'hF3DD] = 8'hC0;
mem[16'hF3DE] = 8'hA9;
mem[16'hF3DF] = 8'h40;
mem[16'hF3E0] = 8'hD0;
mem[16'hF3E1] = 8'h08;
mem[16'hF3E2] = 8'hA9;
mem[16'hF3E3] = 8'h20;
mem[16'hF3E4] = 8'h2C;
mem[16'hF3E5] = 8'h54;
mem[16'hF3E6] = 8'hC0;
mem[16'hF3E7] = 8'h2C;
mem[16'hF3E8] = 8'h53;
mem[16'hF3E9] = 8'hC0;
mem[16'hF3EA] = 8'h85;
mem[16'hF3EB] = 8'hE6;
mem[16'hF3EC] = 8'hAD;
mem[16'hF3ED] = 8'h57;
mem[16'hF3EE] = 8'hC0;
mem[16'hF3EF] = 8'hAD;
mem[16'hF3F0] = 8'h50;
mem[16'hF3F1] = 8'hC0;
mem[16'hF3F2] = 8'hA9;
mem[16'hF3F3] = 8'h00;
mem[16'hF3F4] = 8'h85;
mem[16'hF3F5] = 8'h1C;
mem[16'hF3F6] = 8'hA5;
mem[16'hF3F7] = 8'hE6;
mem[16'hF3F8] = 8'h85;
mem[16'hF3F9] = 8'h1B;
mem[16'hF3FA] = 8'hA0;
mem[16'hF3FB] = 8'h00;
mem[16'hF3FC] = 8'h84;
mem[16'hF3FD] = 8'h1A;
mem[16'hF3FE] = 8'hA5;
mem[16'hF3FF] = 8'h1C;
mem[16'hF400] = 8'h91;
mem[16'hF401] = 8'h1A;
mem[16'hF402] = 8'h20;
mem[16'hF403] = 8'h7E;
mem[16'hF404] = 8'hF4;
mem[16'hF405] = 8'hC8;
mem[16'hF406] = 8'hD0;
mem[16'hF407] = 8'hF6;
mem[16'hF408] = 8'hE6;
mem[16'hF409] = 8'h1B;
mem[16'hF40A] = 8'hA5;
mem[16'hF40B] = 8'h1B;
mem[16'hF40C] = 8'h29;
mem[16'hF40D] = 8'h1F;
mem[16'hF40E] = 8'hD0;
mem[16'hF40F] = 8'hEE;
mem[16'hF410] = 8'h60;
mem[16'hF411] = 8'h85;
mem[16'hF412] = 8'hE2;
mem[16'hF413] = 8'h86;
mem[16'hF414] = 8'hE0;
mem[16'hF415] = 8'h84;
mem[16'hF416] = 8'hE1;
mem[16'hF417] = 8'h48;
mem[16'hF418] = 8'h29;
mem[16'hF419] = 8'hC0;
mem[16'hF41A] = 8'h85;
mem[16'hF41B] = 8'h26;
mem[16'hF41C] = 8'h4A;
mem[16'hF41D] = 8'h4A;
mem[16'hF41E] = 8'h05;
mem[16'hF41F] = 8'h26;
mem[16'hF420] = 8'h85;
mem[16'hF421] = 8'h26;
mem[16'hF422] = 8'h68;
mem[16'hF423] = 8'h85;
mem[16'hF424] = 8'h27;
mem[16'hF425] = 8'h0A;
mem[16'hF426] = 8'h0A;
mem[16'hF427] = 8'h0A;
mem[16'hF428] = 8'h26;
mem[16'hF429] = 8'h27;
mem[16'hF42A] = 8'h0A;
mem[16'hF42B] = 8'h26;
mem[16'hF42C] = 8'h27;
mem[16'hF42D] = 8'h0A;
mem[16'hF42E] = 8'h66;
mem[16'hF42F] = 8'h26;
mem[16'hF430] = 8'hA5;
mem[16'hF431] = 8'h27;
mem[16'hF432] = 8'h29;
mem[16'hF433] = 8'h1F;
mem[16'hF434] = 8'h05;
mem[16'hF435] = 8'hE6;
mem[16'hF436] = 8'h85;
mem[16'hF437] = 8'h27;
mem[16'hF438] = 8'h8A;
mem[16'hF439] = 8'hC0;
mem[16'hF43A] = 8'h00;
mem[16'hF43B] = 8'hF0;
mem[16'hF43C] = 8'h05;
mem[16'hF43D] = 8'hA0;
mem[16'hF43E] = 8'h23;
mem[16'hF43F] = 8'h69;
mem[16'hF440] = 8'h04;
mem[16'hF441] = 8'hC8;
mem[16'hF442] = 8'hE9;
mem[16'hF443] = 8'h07;
mem[16'hF444] = 8'hB0;
mem[16'hF445] = 8'hFB;
mem[16'hF446] = 8'h84;
mem[16'hF447] = 8'hE5;
mem[16'hF448] = 8'hAA;
mem[16'hF449] = 8'hBD;
mem[16'hF44A] = 8'hB9;
mem[16'hF44B] = 8'hF4;
mem[16'hF44C] = 8'h85;
mem[16'hF44D] = 8'h30;
mem[16'hF44E] = 8'h98;
mem[16'hF44F] = 8'h4A;
mem[16'hF450] = 8'hA5;
mem[16'hF451] = 8'hE4;
mem[16'hF452] = 8'h85;
mem[16'hF453] = 8'h1C;
mem[16'hF454] = 8'hB0;
mem[16'hF455] = 8'h28;
mem[16'hF456] = 8'h60;
mem[16'hF457] = 8'h20;
mem[16'hF458] = 8'h11;
mem[16'hF459] = 8'hF4;
mem[16'hF45A] = 8'hA5;
mem[16'hF45B] = 8'h1C;
mem[16'hF45C] = 8'h51;
mem[16'hF45D] = 8'h26;
mem[16'hF45E] = 8'h25;
mem[16'hF45F] = 8'h30;
mem[16'hF460] = 8'h51;
mem[16'hF461] = 8'h26;
mem[16'hF462] = 8'h91;
mem[16'hF463] = 8'h26;
mem[16'hF464] = 8'h60;
mem[16'hF465] = 8'h10;
mem[16'hF466] = 8'h23;
mem[16'hF467] = 8'hA5;
mem[16'hF468] = 8'h30;
mem[16'hF469] = 8'h4A;
mem[16'hF46A] = 8'hB0;
mem[16'hF46B] = 8'h05;
mem[16'hF46C] = 8'h49;
mem[16'hF46D] = 8'hC0;
mem[16'hF46E] = 8'h85;
mem[16'hF46F] = 8'h30;
mem[16'hF470] = 8'h60;
mem[16'hF471] = 8'h88;
mem[16'hF472] = 8'h10;
mem[16'hF473] = 8'h02;
mem[16'hF474] = 8'hA0;
mem[16'hF475] = 8'h27;
mem[16'hF476] = 8'hA9;
mem[16'hF477] = 8'hC0;
mem[16'hF478] = 8'h85;
mem[16'hF479] = 8'h30;
mem[16'hF47A] = 8'h84;
mem[16'hF47B] = 8'hE5;
mem[16'hF47C] = 8'hA5;
mem[16'hF47D] = 8'h1C;
mem[16'hF47E] = 8'h0A;
mem[16'hF47F] = 8'hC9;
mem[16'hF480] = 8'hC0;
mem[16'hF481] = 8'h10;
mem[16'hF482] = 8'h06;
mem[16'hF483] = 8'hA5;
mem[16'hF484] = 8'h1C;
mem[16'hF485] = 8'h49;
mem[16'hF486] = 8'h7F;
mem[16'hF487] = 8'h85;
mem[16'hF488] = 8'h1C;
mem[16'hF489] = 8'h60;
mem[16'hF48A] = 8'hA5;
mem[16'hF48B] = 8'h30;
mem[16'hF48C] = 8'h0A;
mem[16'hF48D] = 8'h49;
mem[16'hF48E] = 8'h80;
mem[16'hF48F] = 8'h30;
mem[16'hF490] = 8'hDD;
mem[16'hF491] = 8'hA9;
mem[16'hF492] = 8'h81;
mem[16'hF493] = 8'hC8;
mem[16'hF494] = 8'hC0;
mem[16'hF495] = 8'h28;
mem[16'hF496] = 8'h90;
mem[16'hF497] = 8'hE0;
mem[16'hF498] = 8'hA0;
mem[16'hF499] = 8'h00;
mem[16'hF49A] = 8'hB0;
mem[16'hF49B] = 8'hDC;
mem[16'hF49C] = 8'h18;
mem[16'hF49D] = 8'hA5;
mem[16'hF49E] = 8'hD1;
mem[16'hF49F] = 8'h29;
mem[16'hF4A0] = 8'h04;
mem[16'hF4A1] = 8'hF0;
mem[16'hF4A2] = 8'h25;
mem[16'hF4A3] = 8'hA9;
mem[16'hF4A4] = 8'h7F;
mem[16'hF4A5] = 8'h25;
mem[16'hF4A6] = 8'h30;
mem[16'hF4A7] = 8'h31;
mem[16'hF4A8] = 8'h26;
mem[16'hF4A9] = 8'hD0;
mem[16'hF4AA] = 8'h19;
mem[16'hF4AB] = 8'hE6;
mem[16'hF4AC] = 8'hEA;
mem[16'hF4AD] = 8'hA9;
mem[16'hF4AE] = 8'h7F;
mem[16'hF4AF] = 8'h25;
mem[16'hF4B0] = 8'h30;
mem[16'hF4B1] = 8'h10;
mem[16'hF4B2] = 8'h11;
mem[16'hF4B3] = 8'h18;
mem[16'hF4B4] = 8'hA5;
mem[16'hF4B5] = 8'hD1;
mem[16'hF4B6] = 8'h29;
mem[16'hF4B7] = 8'h04;
mem[16'hF4B8] = 8'hF0;
mem[16'hF4B9] = 8'h0E;
mem[16'hF4BA] = 8'hB1;
mem[16'hF4BB] = 8'h26;
mem[16'hF4BC] = 8'h45;
mem[16'hF4BD] = 8'h1C;
mem[16'hF4BE] = 8'h25;
mem[16'hF4BF] = 8'h30;
mem[16'hF4C0] = 8'hD0;
mem[16'hF4C1] = 8'h02;
mem[16'hF4C2] = 8'hE6;
mem[16'hF4C3] = 8'hEA;
mem[16'hF4C4] = 8'h51;
mem[16'hF4C5] = 8'h26;
mem[16'hF4C6] = 8'h91;
mem[16'hF4C7] = 8'h26;
mem[16'hF4C8] = 8'hA5;
mem[16'hF4C9] = 8'hD1;
mem[16'hF4CA] = 8'h65;
mem[16'hF4CB] = 8'hD3;
mem[16'hF4CC] = 8'h29;
mem[16'hF4CD] = 8'h03;
mem[16'hF4CE] = 8'hC9;
mem[16'hF4CF] = 8'h02;
mem[16'hF4D0] = 8'h6A;
mem[16'hF4D1] = 8'hB0;
mem[16'hF4D2] = 8'h92;
mem[16'hF4D3] = 8'h30;
mem[16'hF4D4] = 8'h30;
mem[16'hF4D5] = 8'h18;
mem[16'hF4D6] = 8'hA5;
mem[16'hF4D7] = 8'h27;
mem[16'hF4D8] = 8'h2C;
mem[16'hF4D9] = 8'hB9;
mem[16'hF4DA] = 8'hF5;
mem[16'hF4DB] = 8'hD0;
mem[16'hF4DC] = 8'h22;
mem[16'hF4DD] = 8'h06;
mem[16'hF4DE] = 8'h26;
mem[16'hF4DF] = 8'hB0;
mem[16'hF4E0] = 8'h1A;
mem[16'hF4E1] = 8'h2C;
mem[16'hF4E2] = 8'hCD;
mem[16'hF4E3] = 8'hF4;
mem[16'hF4E4] = 8'hF0;
mem[16'hF4E5] = 8'h05;
mem[16'hF4E6] = 8'h69;
mem[16'hF4E7] = 8'h1F;
mem[16'hF4E8] = 8'h38;
mem[16'hF4E9] = 8'hB0;
mem[16'hF4EA] = 8'h12;
mem[16'hF4EB] = 8'h69;
mem[16'hF4EC] = 8'h23;
mem[16'hF4ED] = 8'h48;
mem[16'hF4EE] = 8'hA5;
mem[16'hF4EF] = 8'h26;
mem[16'hF4F0] = 8'h69;
mem[16'hF4F1] = 8'hB0;
mem[16'hF4F2] = 8'hB0;
mem[16'hF4F3] = 8'h02;
mem[16'hF4F4] = 8'h69;
mem[16'hF4F5] = 8'hF0;
mem[16'hF4F6] = 8'h85;
mem[16'hF4F7] = 8'h26;
mem[16'hF4F8] = 8'h68;
mem[16'hF4F9] = 8'hB0;
mem[16'hF4FA] = 8'h02;
mem[16'hF4FB] = 8'h69;
mem[16'hF4FC] = 8'h1F;
mem[16'hF4FD] = 8'h66;
mem[16'hF4FE] = 8'h26;
mem[16'hF4FF] = 8'h69;
mem[16'hF500] = 8'hFC;
mem[16'hF501] = 8'h85;
mem[16'hF502] = 8'h27;
mem[16'hF503] = 8'h60;
mem[16'hF504] = 8'h18;
mem[16'hF505] = 8'hA5;
mem[16'hF506] = 8'h27;
mem[16'hF507] = 8'h69;
mem[16'hF508] = 8'h04;
mem[16'hF509] = 8'h2C;
mem[16'hF50A] = 8'hB9;
mem[16'hF50B] = 8'hF5;
mem[16'hF50C] = 8'hD0;
mem[16'hF50D] = 8'hF3;
mem[16'hF50E] = 8'h06;
mem[16'hF50F] = 8'h26;
mem[16'hF510] = 8'h90;
mem[16'hF511] = 8'h18;
mem[16'hF512] = 8'h69;
mem[16'hF513] = 8'hE0;
mem[16'hF514] = 8'h18;
mem[16'hF515] = 8'h2C;
mem[16'hF516] = 8'h08;
mem[16'hF517] = 8'hF5;
mem[16'hF518] = 8'hF0;
mem[16'hF519] = 8'h12;
mem[16'hF51A] = 8'hA5;
mem[16'hF51B] = 8'h26;
mem[16'hF51C] = 8'h69;
mem[16'hF51D] = 8'h50;
mem[16'hF51E] = 8'h49;
mem[16'hF51F] = 8'hF0;
mem[16'hF520] = 8'hF0;
mem[16'hF521] = 8'h02;
mem[16'hF522] = 8'h49;
mem[16'hF523] = 8'hF0;
mem[16'hF524] = 8'h85;
mem[16'hF525] = 8'h26;
mem[16'hF526] = 8'hA5;
mem[16'hF527] = 8'hE6;
mem[16'hF528] = 8'h90;
mem[16'hF529] = 8'h02;
mem[16'hF52A] = 8'h69;
mem[16'hF52B] = 8'hE0;
mem[16'hF52C] = 8'h66;
mem[16'hF52D] = 8'h26;
mem[16'hF52E] = 8'h90;
mem[16'hF52F] = 8'hD1;
mem[16'hF530] = 8'h48;
mem[16'hF531] = 8'hA9;
mem[16'hF532] = 8'h00;
mem[16'hF533] = 8'h85;
mem[16'hF534] = 8'hE0;
mem[16'hF535] = 8'h85;
mem[16'hF536] = 8'hE1;
mem[16'hF537] = 8'h85;
mem[16'hF538] = 8'hE2;
mem[16'hF539] = 8'h68;
mem[16'hF53A] = 8'h48;
mem[16'hF53B] = 8'h38;
mem[16'hF53C] = 8'hE5;
mem[16'hF53D] = 8'hE0;
mem[16'hF53E] = 8'h48;
mem[16'hF53F] = 8'h8A;
mem[16'hF540] = 8'hE5;
mem[16'hF541] = 8'hE1;
mem[16'hF542] = 8'h85;
mem[16'hF543] = 8'hD3;
mem[16'hF544] = 8'hB0;
mem[16'hF545] = 8'h0A;
mem[16'hF546] = 8'h68;
mem[16'hF547] = 8'h49;
mem[16'hF548] = 8'hFF;
mem[16'hF549] = 8'h69;
mem[16'hF54A] = 8'h01;
mem[16'hF54B] = 8'h48;
mem[16'hF54C] = 8'hA9;
mem[16'hF54D] = 8'h00;
mem[16'hF54E] = 8'hE5;
mem[16'hF54F] = 8'hD3;
mem[16'hF550] = 8'h85;
mem[16'hF551] = 8'hD1;
mem[16'hF552] = 8'h85;
mem[16'hF553] = 8'hD5;
mem[16'hF554] = 8'h68;
mem[16'hF555] = 8'h85;
mem[16'hF556] = 8'hD0;
mem[16'hF557] = 8'h85;
mem[16'hF558] = 8'hD4;
mem[16'hF559] = 8'h68;
mem[16'hF55A] = 8'h85;
mem[16'hF55B] = 8'hE0;
mem[16'hF55C] = 8'h86;
mem[16'hF55D] = 8'hE1;
mem[16'hF55E] = 8'h98;
mem[16'hF55F] = 8'h18;
mem[16'hF560] = 8'hE5;
mem[16'hF561] = 8'hE2;
mem[16'hF562] = 8'h90;
mem[16'hF563] = 8'h04;
mem[16'hF564] = 8'h49;
mem[16'hF565] = 8'hFF;
mem[16'hF566] = 8'h69;
mem[16'hF567] = 8'hFE;
mem[16'hF568] = 8'h85;
mem[16'hF569] = 8'hD2;
mem[16'hF56A] = 8'h84;
mem[16'hF56B] = 8'hE2;
mem[16'hF56C] = 8'h66;
mem[16'hF56D] = 8'hD3;
mem[16'hF56E] = 8'h38;
mem[16'hF56F] = 8'hE5;
mem[16'hF570] = 8'hD0;
mem[16'hF571] = 8'hAA;
mem[16'hF572] = 8'hA9;
mem[16'hF573] = 8'hFF;
mem[16'hF574] = 8'hE5;
mem[16'hF575] = 8'hD1;
mem[16'hF576] = 8'h85;
mem[16'hF577] = 8'h1D;
mem[16'hF578] = 8'hA4;
mem[16'hF579] = 8'hE5;
mem[16'hF57A] = 8'hB0;
mem[16'hF57B] = 8'h05;
mem[16'hF57C] = 8'h0A;
mem[16'hF57D] = 8'h20;
mem[16'hF57E] = 8'h65;
mem[16'hF57F] = 8'hF4;
mem[16'hF580] = 8'h38;
mem[16'hF581] = 8'hA5;
mem[16'hF582] = 8'hD4;
mem[16'hF583] = 8'h65;
mem[16'hF584] = 8'hD2;
mem[16'hF585] = 8'h85;
mem[16'hF586] = 8'hD4;
mem[16'hF587] = 8'hA5;
mem[16'hF588] = 8'hD5;
mem[16'hF589] = 8'hE9;
mem[16'hF58A] = 8'h00;
mem[16'hF58B] = 8'h85;
mem[16'hF58C] = 8'hD5;
mem[16'hF58D] = 8'hB1;
mem[16'hF58E] = 8'h26;
mem[16'hF58F] = 8'h45;
mem[16'hF590] = 8'h1C;
mem[16'hF591] = 8'h25;
mem[16'hF592] = 8'h30;
mem[16'hF593] = 8'h51;
mem[16'hF594] = 8'h26;
mem[16'hF595] = 8'h91;
mem[16'hF596] = 8'h26;
mem[16'hF597] = 8'hE8;
mem[16'hF598] = 8'hD0;
mem[16'hF599] = 8'h04;
mem[16'hF59A] = 8'hE6;
mem[16'hF59B] = 8'h1D;
mem[16'hF59C] = 8'hF0;
mem[16'hF59D] = 8'h62;
mem[16'hF59E] = 8'hA5;
mem[16'hF59F] = 8'hD3;
mem[16'hF5A0] = 8'hB0;
mem[16'hF5A1] = 8'hDA;
mem[16'hF5A2] = 8'h20;
mem[16'hF5A3] = 8'hD3;
mem[16'hF5A4] = 8'hF4;
mem[16'hF5A5] = 8'h18;
mem[16'hF5A6] = 8'hA5;
mem[16'hF5A7] = 8'hD4;
mem[16'hF5A8] = 8'h65;
mem[16'hF5A9] = 8'hD0;
mem[16'hF5AA] = 8'h85;
mem[16'hF5AB] = 8'hD4;
mem[16'hF5AC] = 8'hA5;
mem[16'hF5AD] = 8'hD5;
mem[16'hF5AE] = 8'h65;
mem[16'hF5AF] = 8'hD1;
mem[16'hF5B0] = 8'h50;
mem[16'hF5B1] = 8'hD9;
mem[16'hF5B2] = 8'h81;
mem[16'hF5B3] = 8'h82;
mem[16'hF5B4] = 8'h84;
mem[16'hF5B5] = 8'h88;
mem[16'hF5B6] = 8'h90;
mem[16'hF5B7] = 8'hA0;
mem[16'hF5B8] = 8'hC0;
mem[16'hF5B9] = 8'h1C;
mem[16'hF5BA] = 8'hFF;
mem[16'hF5BB] = 8'hFE;
mem[16'hF5BC] = 8'hFA;
mem[16'hF5BD] = 8'hF4;
mem[16'hF5BE] = 8'hEC;
mem[16'hF5BF] = 8'hE1;
mem[16'hF5C0] = 8'hD4;
mem[16'hF5C1] = 8'hC5;
mem[16'hF5C2] = 8'hB4;
mem[16'hF5C3] = 8'hA1;
mem[16'hF5C4] = 8'h8D;
mem[16'hF5C5] = 8'h78;
mem[16'hF5C6] = 8'h61;
mem[16'hF5C7] = 8'h49;
mem[16'hF5C8] = 8'h31;
mem[16'hF5C9] = 8'h18;
mem[16'hF5CA] = 8'hFF;
mem[16'hF5CB] = 8'hA5;
mem[16'hF5CC] = 8'h26;
mem[16'hF5CD] = 8'h0A;
mem[16'hF5CE] = 8'hA5;
mem[16'hF5CF] = 8'h27;
mem[16'hF5D0] = 8'h29;
mem[16'hF5D1] = 8'h03;
mem[16'hF5D2] = 8'h2A;
mem[16'hF5D3] = 8'h05;
mem[16'hF5D4] = 8'h26;
mem[16'hF5D5] = 8'h0A;
mem[16'hF5D6] = 8'h0A;
mem[16'hF5D7] = 8'h0A;
mem[16'hF5D8] = 8'h85;
mem[16'hF5D9] = 8'hE2;
mem[16'hF5DA] = 8'hA5;
mem[16'hF5DB] = 8'h27;
mem[16'hF5DC] = 8'h4A;
mem[16'hF5DD] = 8'h4A;
mem[16'hF5DE] = 8'h29;
mem[16'hF5DF] = 8'h07;
mem[16'hF5E0] = 8'h05;
mem[16'hF5E1] = 8'hE2;
mem[16'hF5E2] = 8'h85;
mem[16'hF5E3] = 8'hE2;
mem[16'hF5E4] = 8'hA5;
mem[16'hF5E5] = 8'hE5;
mem[16'hF5E6] = 8'h0A;
mem[16'hF5E7] = 8'h65;
mem[16'hF5E8] = 8'hE5;
mem[16'hF5E9] = 8'h0A;
mem[16'hF5EA] = 8'hAA;
mem[16'hF5EB] = 8'hCA;
mem[16'hF5EC] = 8'hA5;
mem[16'hF5ED] = 8'h30;
mem[16'hF5EE] = 8'h29;
mem[16'hF5EF] = 8'h7F;
mem[16'hF5F0] = 8'hE8;
mem[16'hF5F1] = 8'h4A;
mem[16'hF5F2] = 8'hD0;
mem[16'hF5F3] = 8'hFC;
mem[16'hF5F4] = 8'h85;
mem[16'hF5F5] = 8'hE1;
mem[16'hF5F6] = 8'h8A;
mem[16'hF5F7] = 8'h18;
mem[16'hF5F8] = 8'h65;
mem[16'hF5F9] = 8'hE5;
mem[16'hF5FA] = 8'h90;
mem[16'hF5FB] = 8'h02;
mem[16'hF5FC] = 8'hE6;
mem[16'hF5FD] = 8'hE1;
mem[16'hF5FE] = 8'h85;
mem[16'hF5FF] = 8'hE0;
mem[16'hF600] = 8'h60;
mem[16'hF601] = 8'h86;
mem[16'hF602] = 8'h1A;
mem[16'hF603] = 8'h84;
mem[16'hF604] = 8'h1B;
mem[16'hF605] = 8'hAA;
mem[16'hF606] = 8'h4A;
mem[16'hF607] = 8'h4A;
mem[16'hF608] = 8'h4A;
mem[16'hF609] = 8'h4A;
mem[16'hF60A] = 8'h85;
mem[16'hF60B] = 8'hD3;
mem[16'hF60C] = 8'h8A;
mem[16'hF60D] = 8'h29;
mem[16'hF60E] = 8'h0F;
mem[16'hF60F] = 8'hAA;
mem[16'hF610] = 8'hBC;
mem[16'hF611] = 8'hBA;
mem[16'hF612] = 8'hF5;
mem[16'hF613] = 8'h84;
mem[16'hF614] = 8'hD0;
mem[16'hF615] = 8'h49;
mem[16'hF616] = 8'h0F;
mem[16'hF617] = 8'hAA;
mem[16'hF618] = 8'hBC;
mem[16'hF619] = 8'hBB;
mem[16'hF61A] = 8'hF5;
mem[16'hF61B] = 8'hC8;
mem[16'hF61C] = 8'h84;
mem[16'hF61D] = 8'hD2;
mem[16'hF61E] = 8'hA4;
mem[16'hF61F] = 8'hE5;
mem[16'hF620] = 8'hA2;
mem[16'hF621] = 8'h00;
mem[16'hF622] = 8'h86;
mem[16'hF623] = 8'hEA;
mem[16'hF624] = 8'hA1;
mem[16'hF625] = 8'h1A;
mem[16'hF626] = 8'h85;
mem[16'hF627] = 8'hD1;
mem[16'hF628] = 8'hA2;
mem[16'hF629] = 8'h80;
mem[16'hF62A] = 8'h86;
mem[16'hF62B] = 8'hD4;
mem[16'hF62C] = 8'h86;
mem[16'hF62D] = 8'hD5;
mem[16'hF62E] = 8'hA6;
mem[16'hF62F] = 8'hE7;
mem[16'hF630] = 8'hA5;
mem[16'hF631] = 8'hD4;
mem[16'hF632] = 8'h38;
mem[16'hF633] = 8'h65;
mem[16'hF634] = 8'hD0;
mem[16'hF635] = 8'h85;
mem[16'hF636] = 8'hD4;
mem[16'hF637] = 8'h90;
mem[16'hF638] = 8'h04;
mem[16'hF639] = 8'h20;
mem[16'hF63A] = 8'hB3;
mem[16'hF63B] = 8'hF4;
mem[16'hF63C] = 8'h18;
mem[16'hF63D] = 8'hA5;
mem[16'hF63E] = 8'hD5;
mem[16'hF63F] = 8'h65;
mem[16'hF640] = 8'hD2;
mem[16'hF641] = 8'h85;
mem[16'hF642] = 8'hD5;
mem[16'hF643] = 8'h90;
mem[16'hF644] = 8'h03;
mem[16'hF645] = 8'h20;
mem[16'hF646] = 8'hB4;
mem[16'hF647] = 8'hF4;
mem[16'hF648] = 8'hCA;
mem[16'hF649] = 8'hD0;
mem[16'hF64A] = 8'hE5;
mem[16'hF64B] = 8'hA5;
mem[16'hF64C] = 8'hD1;
mem[16'hF64D] = 8'h4A;
mem[16'hF64E] = 8'h4A;
mem[16'hF64F] = 8'h4A;
mem[16'hF650] = 8'hD0;
mem[16'hF651] = 8'hD4;
mem[16'hF652] = 8'hE6;
mem[16'hF653] = 8'h1A;
mem[16'hF654] = 8'hD0;
mem[16'hF655] = 8'h02;
mem[16'hF656] = 8'hE6;
mem[16'hF657] = 8'h1B;
mem[16'hF658] = 8'hA1;
mem[16'hF659] = 8'h1A;
mem[16'hF65A] = 8'hD0;
mem[16'hF65B] = 8'hCA;
mem[16'hF65C] = 8'h60;
mem[16'hF65D] = 8'h86;
mem[16'hF65E] = 8'h1A;
mem[16'hF65F] = 8'h84;
mem[16'hF660] = 8'h1B;
mem[16'hF661] = 8'hAA;
mem[16'hF662] = 8'h4A;
mem[16'hF663] = 8'h4A;
mem[16'hF664] = 8'h4A;
mem[16'hF665] = 8'h4A;
mem[16'hF666] = 8'h85;
mem[16'hF667] = 8'hD3;
mem[16'hF668] = 8'h8A;
mem[16'hF669] = 8'h29;
mem[16'hF66A] = 8'h0F;
mem[16'hF66B] = 8'hAA;
mem[16'hF66C] = 8'hBC;
mem[16'hF66D] = 8'hBA;
mem[16'hF66E] = 8'hF5;
mem[16'hF66F] = 8'h84;
mem[16'hF670] = 8'hD0;
mem[16'hF671] = 8'h49;
mem[16'hF672] = 8'h0F;
mem[16'hF673] = 8'hAA;
mem[16'hF674] = 8'hBC;
mem[16'hF675] = 8'hBB;
mem[16'hF676] = 8'hF5;
mem[16'hF677] = 8'hC8;
mem[16'hF678] = 8'h84;
mem[16'hF679] = 8'hD2;
mem[16'hF67A] = 8'hA4;
mem[16'hF67B] = 8'hE5;
mem[16'hF67C] = 8'hA2;
mem[16'hF67D] = 8'h00;
mem[16'hF67E] = 8'h86;
mem[16'hF67F] = 8'hEA;
mem[16'hF680] = 8'hA1;
mem[16'hF681] = 8'h1A;
mem[16'hF682] = 8'h85;
mem[16'hF683] = 8'hD1;
mem[16'hF684] = 8'hA2;
mem[16'hF685] = 8'h80;
mem[16'hF686] = 8'h86;
mem[16'hF687] = 8'hD4;
mem[16'hF688] = 8'h86;
mem[16'hF689] = 8'hD5;
mem[16'hF68A] = 8'hA6;
mem[16'hF68B] = 8'hE7;
mem[16'hF68C] = 8'hA5;
mem[16'hF68D] = 8'hD4;
mem[16'hF68E] = 8'h38;
mem[16'hF68F] = 8'h65;
mem[16'hF690] = 8'hD0;
mem[16'hF691] = 8'h85;
mem[16'hF692] = 8'hD4;
mem[16'hF693] = 8'h90;
mem[16'hF694] = 8'h04;
mem[16'hF695] = 8'h20;
mem[16'hF696] = 8'h9C;
mem[16'hF697] = 8'hF4;
mem[16'hF698] = 8'h18;
mem[16'hF699] = 8'hA5;
mem[16'hF69A] = 8'hD5;
mem[16'hF69B] = 8'h65;
mem[16'hF69C] = 8'hD2;
mem[16'hF69D] = 8'h85;
mem[16'hF69E] = 8'hD5;
mem[16'hF69F] = 8'h90;
mem[16'hF6A0] = 8'h03;
mem[16'hF6A1] = 8'h20;
mem[16'hF6A2] = 8'h9D;
mem[16'hF6A3] = 8'hF4;
mem[16'hF6A4] = 8'hCA;
mem[16'hF6A5] = 8'hD0;
mem[16'hF6A6] = 8'hE5;
mem[16'hF6A7] = 8'hA5;
mem[16'hF6A8] = 8'hD1;
mem[16'hF6A9] = 8'h4A;
mem[16'hF6AA] = 8'h4A;
mem[16'hF6AB] = 8'h4A;
mem[16'hF6AC] = 8'hD0;
mem[16'hF6AD] = 8'hD4;
mem[16'hF6AE] = 8'hE6;
mem[16'hF6AF] = 8'h1A;
mem[16'hF6B0] = 8'hD0;
mem[16'hF6B1] = 8'h02;
mem[16'hF6B2] = 8'hE6;
mem[16'hF6B3] = 8'h1B;
mem[16'hF6B4] = 8'hA1;
mem[16'hF6B5] = 8'h1A;
mem[16'hF6B6] = 8'hD0;
mem[16'hF6B7] = 8'hCA;
mem[16'hF6B8] = 8'h60;
mem[16'hF6B9] = 8'h20;
mem[16'hF6BA] = 8'h67;
mem[16'hF6BB] = 8'hDD;
mem[16'hF6BC] = 8'h20;
mem[16'hF6BD] = 8'h52;
mem[16'hF6BE] = 8'hE7;
mem[16'hF6BF] = 8'hA4;
mem[16'hF6C0] = 8'h51;
mem[16'hF6C1] = 8'hA6;
mem[16'hF6C2] = 8'h50;
mem[16'hF6C3] = 8'hC0;
mem[16'hF6C4] = 8'h01;
mem[16'hF6C5] = 8'h90;
mem[16'hF6C6] = 8'h06;
mem[16'hF6C7] = 8'hD0;
mem[16'hF6C8] = 8'h1D;
mem[16'hF6C9] = 8'hE0;
mem[16'hF6CA] = 8'h18;
mem[16'hF6CB] = 8'hB0;
mem[16'hF6CC] = 8'h19;
mem[16'hF6CD] = 8'h8A;
mem[16'hF6CE] = 8'h48;
mem[16'hF6CF] = 8'h98;
mem[16'hF6D0] = 8'h48;
mem[16'hF6D1] = 8'hA9;
mem[16'hF6D2] = 8'h2C;
mem[16'hF6D3] = 8'h20;
mem[16'hF6D4] = 8'hC0;
mem[16'hF6D5] = 8'hDE;
mem[16'hF6D6] = 8'h20;
mem[16'hF6D7] = 8'hF8;
mem[16'hF6D8] = 8'hE6;
mem[16'hF6D9] = 8'hE0;
mem[16'hF6DA] = 8'hC0;
mem[16'hF6DB] = 8'hB0;
mem[16'hF6DC] = 8'h09;
mem[16'hF6DD] = 8'h86;
mem[16'hF6DE] = 8'h9D;
mem[16'hF6DF] = 8'h68;
mem[16'hF6E0] = 8'hA8;
mem[16'hF6E1] = 8'h68;
mem[16'hF6E2] = 8'hAA;
mem[16'hF6E3] = 8'hA5;
mem[16'hF6E4] = 8'h9D;
mem[16'hF6E5] = 8'h60;
mem[16'hF6E6] = 8'h4C;
mem[16'hF6E7] = 8'h06;
mem[16'hF6E8] = 8'hF2;
mem[16'hF6E9] = 8'h20;
mem[16'hF6EA] = 8'hF8;
mem[16'hF6EB] = 8'hE6;
mem[16'hF6EC] = 8'hE0;
mem[16'hF6ED] = 8'h08;
mem[16'hF6EE] = 8'hB0;
mem[16'hF6EF] = 8'hF6;
mem[16'hF6F0] = 8'hBD;
mem[16'hF6F1] = 8'hF6;
mem[16'hF6F2] = 8'hF6;
mem[16'hF6F3] = 8'h85;
mem[16'hF6F4] = 8'hE4;
mem[16'hF6F5] = 8'h60;
mem[16'hF6F6] = 8'h00;
mem[16'hF6F7] = 8'h2A;
mem[16'hF6F8] = 8'h55;
mem[16'hF6F9] = 8'h7F;
mem[16'hF6FA] = 8'h80;
mem[16'hF6FB] = 8'hAA;
mem[16'hF6FC] = 8'hD5;
mem[16'hF6FD] = 8'hFF;
mem[16'hF6FE] = 8'hC9;
mem[16'hF6FF] = 8'hC1;
mem[16'hF700] = 8'hF0;
mem[16'hF701] = 8'h0D;
mem[16'hF702] = 8'h20;
mem[16'hF703] = 8'hB9;
mem[16'hF704] = 8'hF6;
mem[16'hF705] = 8'h20;
mem[16'hF706] = 8'h57;
mem[16'hF707] = 8'hF4;
mem[16'hF708] = 8'h20;
mem[16'hF709] = 8'hB7;
mem[16'hF70A] = 8'h00;
mem[16'hF70B] = 8'hC9;
mem[16'hF70C] = 8'hC1;
mem[16'hF70D] = 8'hD0;
mem[16'hF70E] = 8'hE6;
mem[16'hF70F] = 8'h20;
mem[16'hF710] = 8'hC0;
mem[16'hF711] = 8'hDE;
mem[16'hF712] = 8'h20;
mem[16'hF713] = 8'hB9;
mem[16'hF714] = 8'hF6;
mem[16'hF715] = 8'h84;
mem[16'hF716] = 8'h9D;
mem[16'hF717] = 8'hA8;
mem[16'hF718] = 8'h8A;
mem[16'hF719] = 8'hA6;
mem[16'hF71A] = 8'h9D;
mem[16'hF71B] = 8'h20;
mem[16'hF71C] = 8'h3A;
mem[16'hF71D] = 8'hF5;
mem[16'hF71E] = 8'h4C;
mem[16'hF71F] = 8'h08;
mem[16'hF720] = 8'hF7;
mem[16'hF721] = 8'h20;
mem[16'hF722] = 8'hF8;
mem[16'hF723] = 8'hE6;
mem[16'hF724] = 8'h86;
mem[16'hF725] = 8'hF9;
mem[16'hF726] = 8'h60;
mem[16'hF727] = 8'h20;
mem[16'hF728] = 8'hF8;
mem[16'hF729] = 8'hE6;
mem[16'hF72A] = 8'h86;
mem[16'hF72B] = 8'hE7;
mem[16'hF72C] = 8'h60;
mem[16'hF72D] = 8'h20;
mem[16'hF72E] = 8'hF8;
mem[16'hF72F] = 8'hE6;
mem[16'hF730] = 8'hA5;
mem[16'hF731] = 8'hE8;
mem[16'hF732] = 8'h85;
mem[16'hF733] = 8'h1A;
mem[16'hF734] = 8'hA5;
mem[16'hF735] = 8'hE9;
mem[16'hF736] = 8'h85;
mem[16'hF737] = 8'h1B;
mem[16'hF738] = 8'h8A;
mem[16'hF739] = 8'hA2;
mem[16'hF73A] = 8'h00;
mem[16'hF73B] = 8'hC1;
mem[16'hF73C] = 8'h1A;
mem[16'hF73D] = 8'hF0;
mem[16'hF73E] = 8'h02;
mem[16'hF73F] = 8'hB0;
mem[16'hF740] = 8'hA5;
mem[16'hF741] = 8'h0A;
mem[16'hF742] = 8'h90;
mem[16'hF743] = 8'h03;
mem[16'hF744] = 8'hE6;
mem[16'hF745] = 8'h1B;
mem[16'hF746] = 8'h18;
mem[16'hF747] = 8'hA8;
mem[16'hF748] = 8'hB1;
mem[16'hF749] = 8'h1A;
mem[16'hF74A] = 8'h65;
mem[16'hF74B] = 8'h1A;
mem[16'hF74C] = 8'hAA;
mem[16'hF74D] = 8'hC8;
mem[16'hF74E] = 8'hB1;
mem[16'hF74F] = 8'h1A;
mem[16'hF750] = 8'h65;
mem[16'hF751] = 8'hE9;
mem[16'hF752] = 8'h85;
mem[16'hF753] = 8'h1B;
mem[16'hF754] = 8'h86;
mem[16'hF755] = 8'h1A;
mem[16'hF756] = 8'h20;
mem[16'hF757] = 8'hB7;
mem[16'hF758] = 8'h00;
mem[16'hF759] = 8'hC9;
mem[16'hF75A] = 8'hC5;
mem[16'hF75B] = 8'hD0;
mem[16'hF75C] = 8'h09;
mem[16'hF75D] = 8'h20;
mem[16'hF75E] = 8'hC0;
mem[16'hF75F] = 8'hDE;
mem[16'hF760] = 8'h20;
mem[16'hF761] = 8'hB9;
mem[16'hF762] = 8'hF6;
mem[16'hF763] = 8'h20;
mem[16'hF764] = 8'h11;
mem[16'hF765] = 8'hF4;
mem[16'hF766] = 8'hA5;
mem[16'hF767] = 8'hF9;
mem[16'hF768] = 8'h60;
mem[16'hF769] = 8'h20;
mem[16'hF76A] = 8'h2D;
mem[16'hF76B] = 8'hF7;
mem[16'hF76C] = 8'h4C;
mem[16'hF76D] = 8'h05;
mem[16'hF76E] = 8'hF6;
mem[16'hF76F] = 8'h20;
mem[16'hF770] = 8'h2D;
mem[16'hF771] = 8'hF7;
mem[16'hF772] = 8'h4C;
mem[16'hF773] = 8'h61;
mem[16'hF774] = 8'hF6;
mem[16'hF775] = 8'hA9;
mem[16'hF776] = 8'h00;
mem[16'hF777] = 8'h85;
mem[16'hF778] = 8'h3D;
mem[16'hF779] = 8'h85;
mem[16'hF77A] = 8'h3F;
mem[16'hF77B] = 8'hA0;
mem[16'hF77C] = 8'h50;
mem[16'hF77D] = 8'h84;
mem[16'hF77E] = 8'h3C;
mem[16'hF77F] = 8'hC8;
mem[16'hF780] = 8'h84;
mem[16'hF781] = 8'h3E;
mem[16'hF782] = 8'h20;
mem[16'hF783] = 8'hFD;
mem[16'hF784] = 8'hFE;
mem[16'hF785] = 8'h18;
mem[16'hF786] = 8'hA5;
mem[16'hF787] = 8'h73;
mem[16'hF788] = 8'hAA;
mem[16'hF789] = 8'hCA;
mem[16'hF78A] = 8'h86;
mem[16'hF78B] = 8'h3E;
mem[16'hF78C] = 8'hE5;
mem[16'hF78D] = 8'h50;
mem[16'hF78E] = 8'h48;
mem[16'hF78F] = 8'hA5;
mem[16'hF790] = 8'h74;
mem[16'hF791] = 8'hA8;
mem[16'hF792] = 8'hE8;
mem[16'hF793] = 8'hD0;
mem[16'hF794] = 8'h01;
mem[16'hF795] = 8'h88;
mem[16'hF796] = 8'h84;
mem[16'hF797] = 8'h3F;
mem[16'hF798] = 8'hE5;
mem[16'hF799] = 8'h51;
mem[16'hF79A] = 8'hC5;
mem[16'hF79B] = 8'h6E;
mem[16'hF79C] = 8'h90;
mem[16'hF79D] = 8'h02;
mem[16'hF79E] = 8'hD0;
mem[16'hF79F] = 8'h03;
mem[16'hF7A0] = 8'h4C;
mem[16'hF7A1] = 8'h10;
mem[16'hF7A2] = 8'hD4;
mem[16'hF7A3] = 8'h85;
mem[16'hF7A4] = 8'h74;
mem[16'hF7A5] = 8'h85;
mem[16'hF7A6] = 8'h70;
mem[16'hF7A7] = 8'h85;
mem[16'hF7A8] = 8'h3D;
mem[16'hF7A9] = 8'h85;
mem[16'hF7AA] = 8'hE9;
mem[16'hF7AB] = 8'h68;
mem[16'hF7AC] = 8'h85;
mem[16'hF7AD] = 8'hE8;
mem[16'hF7AE] = 8'h85;
mem[16'hF7AF] = 8'h73;
mem[16'hF7B0] = 8'h85;
mem[16'hF7B1] = 8'h6F;
mem[16'hF7B2] = 8'h85;
mem[16'hF7B3] = 8'h3C;
mem[16'hF7B4] = 8'h20;
mem[16'hF7B5] = 8'hFA;
mem[16'hF7B6] = 8'hFC;
mem[16'hF7B7] = 8'hA9;
mem[16'hF7B8] = 8'h03;
mem[16'hF7B9] = 8'h4C;
mem[16'hF7BA] = 8'h02;
mem[16'hF7BB] = 8'hFF;
mem[16'hF7BC] = 8'h18;
mem[16'hF7BD] = 8'hA5;
mem[16'hF7BE] = 8'h9B;
mem[16'hF7BF] = 8'h65;
mem[16'hF7C0] = 8'h50;
mem[16'hF7C1] = 8'h85;
mem[16'hF7C2] = 8'h3E;
mem[16'hF7C3] = 8'hA5;
mem[16'hF7C4] = 8'h9C;
mem[16'hF7C5] = 8'h65;
mem[16'hF7C6] = 8'h51;
mem[16'hF7C7] = 8'h85;
mem[16'hF7C8] = 8'h3F;
mem[16'hF7C9] = 8'hA0;
mem[16'hF7CA] = 8'h04;
mem[16'hF7CB] = 8'hB1;
mem[16'hF7CC] = 8'h9B;
mem[16'hF7CD] = 8'h20;
mem[16'hF7CE] = 8'hEF;
mem[16'hF7CF] = 8'hE0;
mem[16'hF7D0] = 8'hA5;
mem[16'hF7D1] = 8'h94;
mem[16'hF7D2] = 8'h85;
mem[16'hF7D3] = 8'h3C;
mem[16'hF7D4] = 8'hA5;
mem[16'hF7D5] = 8'h95;
mem[16'hF7D6] = 8'h85;
mem[16'hF7D7] = 8'h3D;
mem[16'hF7D8] = 8'h60;
mem[16'hF7D9] = 8'hA9;
mem[16'hF7DA] = 8'h40;
mem[16'hF7DB] = 8'h85;
mem[16'hF7DC] = 8'h14;
mem[16'hF7DD] = 8'h20;
mem[16'hF7DE] = 8'hE3;
mem[16'hF7DF] = 8'hDF;
mem[16'hF7E0] = 8'hA9;
mem[16'hF7E1] = 8'h00;
mem[16'hF7E2] = 8'h85;
mem[16'hF7E3] = 8'h14;
mem[16'hF7E4] = 8'h4C;
mem[16'hF7E5] = 8'hF0;
mem[16'hF7E6] = 8'hD8;
mem[16'hF7E7] = 8'h20;
mem[16'hF7E8] = 8'hF8;
mem[16'hF7E9] = 8'hE6;
mem[16'hF7EA] = 8'hCA;
mem[16'hF7EB] = 8'h8A;
mem[16'hF7EC] = 8'hC9;
mem[16'hF7ED] = 8'h28;
mem[16'hF7EE] = 8'h90;
mem[16'hF7EF] = 8'h0A;
mem[16'hF7F0] = 8'hE9;
mem[16'hF7F1] = 8'h28;
mem[16'hF7F2] = 8'h48;
mem[16'hF7F3] = 8'h20;
mem[16'hF7F4] = 8'hFB;
mem[16'hF7F5] = 8'hDA;
mem[16'hF7F6] = 8'h68;
mem[16'hF7F7] = 8'h4C;
mem[16'hF7F8] = 8'hEC;
mem[16'hF7F9] = 8'hF7;
mem[16'hF7FA] = 8'h85;
mem[16'hF7FB] = 8'h24;
mem[16'hF7FC] = 8'h60;
mem[16'hF7FD] = 8'hCB;
mem[16'hF7FE] = 8'hD2;
mem[16'hF7FF] = 8'h78;
mem[16'hF800] = 8'h4A;
mem[16'hF801] = 8'h08;
mem[16'hF802] = 8'h20;
mem[16'hF803] = 8'h47;
mem[16'hF804] = 8'hF8;
mem[16'hF805] = 8'h28;
mem[16'hF806] = 8'hA9;
mem[16'hF807] = 8'h0F;
mem[16'hF808] = 8'h90;
mem[16'hF809] = 8'h02;
mem[16'hF80A] = 8'h69;
mem[16'hF80B] = 8'hE0;
mem[16'hF80C] = 8'h85;
mem[16'hF80D] = 8'h2E;
mem[16'hF80E] = 8'hB1;
mem[16'hF80F] = 8'h26;
mem[16'hF810] = 8'h45;
mem[16'hF811] = 8'h30;
mem[16'hF812] = 8'h25;
mem[16'hF813] = 8'h2E;
mem[16'hF814] = 8'h51;
mem[16'hF815] = 8'h26;
mem[16'hF816] = 8'h91;
mem[16'hF817] = 8'h26;
mem[16'hF818] = 8'h60;
mem[16'hF819] = 8'h20;
mem[16'hF81A] = 8'h00;
mem[16'hF81B] = 8'hF8;
mem[16'hF81C] = 8'hC4;
mem[16'hF81D] = 8'h2C;
mem[16'hF81E] = 8'hB0;
mem[16'hF81F] = 8'h11;
mem[16'hF820] = 8'hC8;
mem[16'hF821] = 8'h20;
mem[16'hF822] = 8'h0E;
mem[16'hF823] = 8'hF8;
mem[16'hF824] = 8'h90;
mem[16'hF825] = 8'hF6;
mem[16'hF826] = 8'h69;
mem[16'hF827] = 8'h01;
mem[16'hF828] = 8'h48;
mem[16'hF829] = 8'h20;
mem[16'hF82A] = 8'h00;
mem[16'hF82B] = 8'hF8;
mem[16'hF82C] = 8'h68;
mem[16'hF82D] = 8'hC5;
mem[16'hF82E] = 8'h2D;
mem[16'hF82F] = 8'h90;
mem[16'hF830] = 8'hF5;
mem[16'hF831] = 8'h60;
mem[16'hF832] = 8'hA0;
mem[16'hF833] = 8'h2F;
mem[16'hF834] = 8'hD0;
mem[16'hF835] = 8'h02;
mem[16'hF836] = 8'hA0;
mem[16'hF837] = 8'h27;
mem[16'hF838] = 8'h84;
mem[16'hF839] = 8'h2D;
mem[16'hF83A] = 8'hA0;
mem[16'hF83B] = 8'h27;
mem[16'hF83C] = 8'hA9;
mem[16'hF83D] = 8'h00;
mem[16'hF83E] = 8'h85;
mem[16'hF83F] = 8'h30;
mem[16'hF840] = 8'h20;
mem[16'hF841] = 8'h28;
mem[16'hF842] = 8'hF8;
mem[16'hF843] = 8'h88;
mem[16'hF844] = 8'h10;
mem[16'hF845] = 8'hF6;
mem[16'hF846] = 8'h60;
mem[16'hF847] = 8'h48;
mem[16'hF848] = 8'h4A;
mem[16'hF849] = 8'h29;
mem[16'hF84A] = 8'h03;
mem[16'hF84B] = 8'h09;
mem[16'hF84C] = 8'h04;
mem[16'hF84D] = 8'h85;
mem[16'hF84E] = 8'h27;
mem[16'hF84F] = 8'h68;
mem[16'hF850] = 8'h29;
mem[16'hF851] = 8'h18;
mem[16'hF852] = 8'h90;
mem[16'hF853] = 8'h02;
mem[16'hF854] = 8'h69;
mem[16'hF855] = 8'h7F;
mem[16'hF856] = 8'h85;
mem[16'hF857] = 8'h26;
mem[16'hF858] = 8'h0A;
mem[16'hF859] = 8'h0A;
mem[16'hF85A] = 8'h05;
mem[16'hF85B] = 8'h26;
mem[16'hF85C] = 8'h85;
mem[16'hF85D] = 8'h26;
mem[16'hF85E] = 8'h60;
mem[16'hF85F] = 8'hA5;
mem[16'hF860] = 8'h30;
mem[16'hF861] = 8'h18;
mem[16'hF862] = 8'h69;
mem[16'hF863] = 8'h03;
mem[16'hF864] = 8'h29;
mem[16'hF865] = 8'h0F;
mem[16'hF866] = 8'h85;
mem[16'hF867] = 8'h30;
mem[16'hF868] = 8'h0A;
mem[16'hF869] = 8'h0A;
mem[16'hF86A] = 8'h0A;
mem[16'hF86B] = 8'h0A;
mem[16'hF86C] = 8'h05;
mem[16'hF86D] = 8'h30;
mem[16'hF86E] = 8'h85;
mem[16'hF86F] = 8'h30;
mem[16'hF870] = 8'h60;
mem[16'hF871] = 8'h4A;
mem[16'hF872] = 8'h08;
mem[16'hF873] = 8'h20;
mem[16'hF874] = 8'h47;
mem[16'hF875] = 8'hF8;
mem[16'hF876] = 8'hB1;
mem[16'hF877] = 8'h26;
mem[16'hF878] = 8'h28;
mem[16'hF879] = 8'h90;
mem[16'hF87A] = 8'h04;
mem[16'hF87B] = 8'h4A;
mem[16'hF87C] = 8'h4A;
mem[16'hF87D] = 8'h4A;
mem[16'hF87E] = 8'h4A;
mem[16'hF87F] = 8'h29;
mem[16'hF880] = 8'h0F;
mem[16'hF881] = 8'h60;
mem[16'hF882] = 8'hA6;
mem[16'hF883] = 8'h3A;
mem[16'hF884] = 8'hA4;
mem[16'hF885] = 8'h3B;
mem[16'hF886] = 8'h20;
mem[16'hF887] = 8'h96;
mem[16'hF888] = 8'hFD;
mem[16'hF889] = 8'h20;
mem[16'hF88A] = 8'h48;
mem[16'hF88B] = 8'hF9;
mem[16'hF88C] = 8'hA1;
mem[16'hF88D] = 8'h3A;
mem[16'hF88E] = 8'hA8;
mem[16'hF88F] = 8'h4A;
mem[16'hF890] = 8'h90;
mem[16'hF891] = 8'h09;
mem[16'hF892] = 8'h6A;
mem[16'hF893] = 8'hB0;
mem[16'hF894] = 8'h10;
mem[16'hF895] = 8'hC9;
mem[16'hF896] = 8'hA2;
mem[16'hF897] = 8'hF0;
mem[16'hF898] = 8'h0C;
mem[16'hF899] = 8'h29;
mem[16'hF89A] = 8'h87;
mem[16'hF89B] = 8'h4A;
mem[16'hF89C] = 8'hAA;
mem[16'hF89D] = 8'hBD;
mem[16'hF89E] = 8'h62;
mem[16'hF89F] = 8'hF9;
mem[16'hF8A0] = 8'h20;
mem[16'hF8A1] = 8'h79;
mem[16'hF8A2] = 8'hF8;
mem[16'hF8A3] = 8'hD0;
mem[16'hF8A4] = 8'h04;
mem[16'hF8A5] = 8'hA0;
mem[16'hF8A6] = 8'h80;
mem[16'hF8A7] = 8'hA9;
mem[16'hF8A8] = 8'h00;
mem[16'hF8A9] = 8'hAA;
mem[16'hF8AA] = 8'hBD;
mem[16'hF8AB] = 8'hA6;
mem[16'hF8AC] = 8'hF9;
mem[16'hF8AD] = 8'h85;
mem[16'hF8AE] = 8'h2E;
mem[16'hF8AF] = 8'h29;
mem[16'hF8B0] = 8'h03;
mem[16'hF8B1] = 8'h85;
mem[16'hF8B2] = 8'h2F;
mem[16'hF8B3] = 8'h98;
mem[16'hF8B4] = 8'h29;
mem[16'hF8B5] = 8'h8F;
mem[16'hF8B6] = 8'hAA;
mem[16'hF8B7] = 8'h98;
mem[16'hF8B8] = 8'hA0;
mem[16'hF8B9] = 8'h03;
mem[16'hF8BA] = 8'hE0;
mem[16'hF8BB] = 8'h8A;
mem[16'hF8BC] = 8'hF0;
mem[16'hF8BD] = 8'h0B;
mem[16'hF8BE] = 8'h4A;
mem[16'hF8BF] = 8'h90;
mem[16'hF8C0] = 8'h08;
mem[16'hF8C1] = 8'h4A;
mem[16'hF8C2] = 8'h4A;
mem[16'hF8C3] = 8'h09;
mem[16'hF8C4] = 8'h20;
mem[16'hF8C5] = 8'h88;
mem[16'hF8C6] = 8'hD0;
mem[16'hF8C7] = 8'hFA;
mem[16'hF8C8] = 8'hC8;
mem[16'hF8C9] = 8'h88;
mem[16'hF8CA] = 8'hD0;
mem[16'hF8CB] = 8'hF2;
mem[16'hF8CC] = 8'h60;
mem[16'hF8CD] = 8'hFF;
mem[16'hF8CE] = 8'hFF;
mem[16'hF8CF] = 8'hFF;
mem[16'hF8D0] = 8'h20;
mem[16'hF8D1] = 8'h82;
mem[16'hF8D2] = 8'hF8;
mem[16'hF8D3] = 8'h48;
mem[16'hF8D4] = 8'hB1;
mem[16'hF8D5] = 8'h3A;
mem[16'hF8D6] = 8'h20;
mem[16'hF8D7] = 8'hDA;
mem[16'hF8D8] = 8'hFD;
mem[16'hF8D9] = 8'hA2;
mem[16'hF8DA] = 8'h01;
mem[16'hF8DB] = 8'h20;
mem[16'hF8DC] = 8'h4A;
mem[16'hF8DD] = 8'hF9;
mem[16'hF8DE] = 8'hC4;
mem[16'hF8DF] = 8'h2F;
mem[16'hF8E0] = 8'hC8;
mem[16'hF8E1] = 8'h90;
mem[16'hF8E2] = 8'hF1;
mem[16'hF8E3] = 8'hA2;
mem[16'hF8E4] = 8'h03;
mem[16'hF8E5] = 8'hC0;
mem[16'hF8E6] = 8'h04;
mem[16'hF8E7] = 8'h90;
mem[16'hF8E8] = 8'hF2;
mem[16'hF8E9] = 8'h68;
mem[16'hF8EA] = 8'hA8;
mem[16'hF8EB] = 8'hB9;
mem[16'hF8EC] = 8'hC0;
mem[16'hF8ED] = 8'hF9;
mem[16'hF8EE] = 8'h85;
mem[16'hF8EF] = 8'h2C;
mem[16'hF8F0] = 8'hB9;
mem[16'hF8F1] = 8'h00;
mem[16'hF8F2] = 8'hFA;
mem[16'hF8F3] = 8'h85;
mem[16'hF8F4] = 8'h2D;
mem[16'hF8F5] = 8'hA9;
mem[16'hF8F6] = 8'h00;
mem[16'hF8F7] = 8'hA0;
mem[16'hF8F8] = 8'h05;
mem[16'hF8F9] = 8'h06;
mem[16'hF8FA] = 8'h2D;
mem[16'hF8FB] = 8'h26;
mem[16'hF8FC] = 8'h2C;
mem[16'hF8FD] = 8'h2A;
mem[16'hF8FE] = 8'h88;
mem[16'hF8FF] = 8'hD0;
mem[16'hF900] = 8'hF8;
mem[16'hF901] = 8'h69;
mem[16'hF902] = 8'hBF;
mem[16'hF903] = 8'h20;
mem[16'hF904] = 8'hED;
mem[16'hF905] = 8'hFD;
mem[16'hF906] = 8'hCA;
mem[16'hF907] = 8'hD0;
mem[16'hF908] = 8'hEC;
mem[16'hF909] = 8'h20;
mem[16'hF90A] = 8'h48;
mem[16'hF90B] = 8'hF9;
mem[16'hF90C] = 8'hA4;
mem[16'hF90D] = 8'h2F;
mem[16'hF90E] = 8'hA2;
mem[16'hF90F] = 8'h06;
mem[16'hF910] = 8'hE0;
mem[16'hF911] = 8'h03;
mem[16'hF912] = 8'hF0;
mem[16'hF913] = 8'h1C;
mem[16'hF914] = 8'h06;
mem[16'hF915] = 8'h2E;
mem[16'hF916] = 8'h90;
mem[16'hF917] = 8'h0E;
mem[16'hF918] = 8'hBD;
mem[16'hF919] = 8'hB3;
mem[16'hF91A] = 8'hF9;
mem[16'hF91B] = 8'h20;
mem[16'hF91C] = 8'hED;
mem[16'hF91D] = 8'hFD;
mem[16'hF91E] = 8'hBD;
mem[16'hF91F] = 8'hB9;
mem[16'hF920] = 8'hF9;
mem[16'hF921] = 8'hF0;
mem[16'hF922] = 8'h03;
mem[16'hF923] = 8'h20;
mem[16'hF924] = 8'hED;
mem[16'hF925] = 8'hFD;
mem[16'hF926] = 8'hCA;
mem[16'hF927] = 8'hD0;
mem[16'hF928] = 8'hE7;
mem[16'hF929] = 8'h60;
mem[16'hF92A] = 8'h88;
mem[16'hF92B] = 8'h30;
mem[16'hF92C] = 8'hE7;
mem[16'hF92D] = 8'h20;
mem[16'hF92E] = 8'hDA;
mem[16'hF92F] = 8'hFD;
mem[16'hF930] = 8'hA5;
mem[16'hF931] = 8'h2E;
mem[16'hF932] = 8'hC9;
mem[16'hF933] = 8'hE8;
mem[16'hF934] = 8'hB1;
mem[16'hF935] = 8'h3A;
mem[16'hF936] = 8'h90;
mem[16'hF937] = 8'hF2;
mem[16'hF938] = 8'h20;
mem[16'hF939] = 8'h56;
mem[16'hF93A] = 8'hF9;
mem[16'hF93B] = 8'hAA;
mem[16'hF93C] = 8'hE8;
mem[16'hF93D] = 8'hD0;
mem[16'hF93E] = 8'h01;
mem[16'hF93F] = 8'hC8;
mem[16'hF940] = 8'h98;
mem[16'hF941] = 8'h20;
mem[16'hF942] = 8'hDA;
mem[16'hF943] = 8'hFD;
mem[16'hF944] = 8'h8A;
mem[16'hF945] = 8'h4C;
mem[16'hF946] = 8'hDA;
mem[16'hF947] = 8'hFD;
mem[16'hF948] = 8'hA2;
mem[16'hF949] = 8'h03;
mem[16'hF94A] = 8'hA9;
mem[16'hF94B] = 8'hA0;
mem[16'hF94C] = 8'h20;
mem[16'hF94D] = 8'hED;
mem[16'hF94E] = 8'hFD;
mem[16'hF94F] = 8'hCA;
mem[16'hF950] = 8'hD0;
mem[16'hF951] = 8'hF8;
mem[16'hF952] = 8'h60;
mem[16'hF953] = 8'h38;
mem[16'hF954] = 8'hA5;
mem[16'hF955] = 8'h2F;
mem[16'hF956] = 8'hA4;
mem[16'hF957] = 8'h3B;
mem[16'hF958] = 8'hAA;
mem[16'hF959] = 8'h10;
mem[16'hF95A] = 8'h01;
mem[16'hF95B] = 8'h88;
mem[16'hF95C] = 8'h65;
mem[16'hF95D] = 8'h3A;
mem[16'hF95E] = 8'h90;
mem[16'hF95F] = 8'h01;
mem[16'hF960] = 8'hC8;
mem[16'hF961] = 8'h60;
mem[16'hF962] = 8'h04;
mem[16'hF963] = 8'h20;
mem[16'hF964] = 8'h54;
mem[16'hF965] = 8'h30;
mem[16'hF966] = 8'h0D;
mem[16'hF967] = 8'h80;
mem[16'hF968] = 8'h04;
mem[16'hF969] = 8'h90;
mem[16'hF96A] = 8'h03;
mem[16'hF96B] = 8'h22;
mem[16'hF96C] = 8'h54;
mem[16'hF96D] = 8'h33;
mem[16'hF96E] = 8'h0D;
mem[16'hF96F] = 8'h80;
mem[16'hF970] = 8'h04;
mem[16'hF971] = 8'h90;
mem[16'hF972] = 8'h04;
mem[16'hF973] = 8'h20;
mem[16'hF974] = 8'h54;
mem[16'hF975] = 8'h33;
mem[16'hF976] = 8'h0D;
mem[16'hF977] = 8'h80;
mem[16'hF978] = 8'h04;
mem[16'hF979] = 8'h90;
mem[16'hF97A] = 8'h04;
mem[16'hF97B] = 8'h20;
mem[16'hF97C] = 8'h54;
mem[16'hF97D] = 8'h3B;
mem[16'hF97E] = 8'h0D;
mem[16'hF97F] = 8'h80;
mem[16'hF980] = 8'h04;
mem[16'hF981] = 8'h90;
mem[16'hF982] = 8'h00;
mem[16'hF983] = 8'h22;
mem[16'hF984] = 8'h44;
mem[16'hF985] = 8'h33;
mem[16'hF986] = 8'h0D;
mem[16'hF987] = 8'hC8;
mem[16'hF988] = 8'h44;
mem[16'hF989] = 8'h00;
mem[16'hF98A] = 8'h11;
mem[16'hF98B] = 8'h22;
mem[16'hF98C] = 8'h44;
mem[16'hF98D] = 8'h33;
mem[16'hF98E] = 8'h0D;
mem[16'hF98F] = 8'hC8;
mem[16'hF990] = 8'h44;
mem[16'hF991] = 8'hA9;
mem[16'hF992] = 8'h01;
mem[16'hF993] = 8'h22;
mem[16'hF994] = 8'h44;
mem[16'hF995] = 8'h33;
mem[16'hF996] = 8'h0D;
mem[16'hF997] = 8'h80;
mem[16'hF998] = 8'h04;
mem[16'hF999] = 8'h90;
mem[16'hF99A] = 8'h01;
mem[16'hF99B] = 8'h22;
mem[16'hF99C] = 8'h44;
mem[16'hF99D] = 8'h33;
mem[16'hF99E] = 8'h0D;
mem[16'hF99F] = 8'h80;
mem[16'hF9A0] = 8'h04;
mem[16'hF9A1] = 8'h90;
mem[16'hF9A2] = 8'h26;
mem[16'hF9A3] = 8'h31;
mem[16'hF9A4] = 8'h87;
mem[16'hF9A5] = 8'h9A;
mem[16'hF9A6] = 8'h00;
mem[16'hF9A7] = 8'h21;
mem[16'hF9A8] = 8'h81;
mem[16'hF9A9] = 8'h82;
mem[16'hF9AA] = 8'h00;
mem[16'hF9AB] = 8'h00;
mem[16'hF9AC] = 8'h59;
mem[16'hF9AD] = 8'h4D;
mem[16'hF9AE] = 8'h91;
mem[16'hF9AF] = 8'h92;
mem[16'hF9B0] = 8'h86;
mem[16'hF9B1] = 8'h4A;
mem[16'hF9B2] = 8'h85;
mem[16'hF9B3] = 8'h9D;
mem[16'hF9B4] = 8'hAC;
mem[16'hF9B5] = 8'hA9;
mem[16'hF9B6] = 8'hAC;
mem[16'hF9B7] = 8'hA3;
mem[16'hF9B8] = 8'hA8;
mem[16'hF9B9] = 8'hA4;
mem[16'hF9BA] = 8'hD9;
mem[16'hF9BB] = 8'h00;
mem[16'hF9BC] = 8'hD8;
mem[16'hF9BD] = 8'hA4;
mem[16'hF9BE] = 8'hA4;
mem[16'hF9BF] = 8'h00;
mem[16'hF9C0] = 8'h1C;
mem[16'hF9C1] = 8'h8A;
mem[16'hF9C2] = 8'h1C;
mem[16'hF9C3] = 8'h23;
mem[16'hF9C4] = 8'h5D;
mem[16'hF9C5] = 8'h8B;
mem[16'hF9C6] = 8'h1B;
mem[16'hF9C7] = 8'hA1;
mem[16'hF9C8] = 8'h9D;
mem[16'hF9C9] = 8'h8A;
mem[16'hF9CA] = 8'h1D;
mem[16'hF9CB] = 8'h23;
mem[16'hF9CC] = 8'h9D;
mem[16'hF9CD] = 8'h8B;
mem[16'hF9CE] = 8'h1D;
mem[16'hF9CF] = 8'hA1;
mem[16'hF9D0] = 8'h00;
mem[16'hF9D1] = 8'h29;
mem[16'hF9D2] = 8'h19;
mem[16'hF9D3] = 8'hAE;
mem[16'hF9D4] = 8'h69;
mem[16'hF9D5] = 8'hA8;
mem[16'hF9D6] = 8'h19;
mem[16'hF9D7] = 8'h23;
mem[16'hF9D8] = 8'h24;
mem[16'hF9D9] = 8'h53;
mem[16'hF9DA] = 8'h1B;
mem[16'hF9DB] = 8'h23;
mem[16'hF9DC] = 8'h24;
mem[16'hF9DD] = 8'h53;
mem[16'hF9DE] = 8'h19;
mem[16'hF9DF] = 8'hA1;
mem[16'hF9E0] = 8'h00;
mem[16'hF9E1] = 8'h1A;
mem[16'hF9E2] = 8'h5B;
mem[16'hF9E3] = 8'h5B;
mem[16'hF9E4] = 8'hA5;
mem[16'hF9E5] = 8'h69;
mem[16'hF9E6] = 8'h24;
mem[16'hF9E7] = 8'h24;
mem[16'hF9E8] = 8'hAE;
mem[16'hF9E9] = 8'hAE;
mem[16'hF9EA] = 8'hA8;
mem[16'hF9EB] = 8'hAD;
mem[16'hF9EC] = 8'h29;
mem[16'hF9ED] = 8'h00;
mem[16'hF9EE] = 8'h7C;
mem[16'hF9EF] = 8'h00;
mem[16'hF9F0] = 8'h15;
mem[16'hF9F1] = 8'h9C;
mem[16'hF9F2] = 8'h6D;
mem[16'hF9F3] = 8'h9C;
mem[16'hF9F4] = 8'hA5;
mem[16'hF9F5] = 8'h69;
mem[16'hF9F6] = 8'h29;
mem[16'hF9F7] = 8'h53;
mem[16'hF9F8] = 8'h84;
mem[16'hF9F9] = 8'h13;
mem[16'hF9FA] = 8'h34;
mem[16'hF9FB] = 8'h11;
mem[16'hF9FC] = 8'hA5;
mem[16'hF9FD] = 8'h69;
mem[16'hF9FE] = 8'h23;
mem[16'hF9FF] = 8'hA0;
mem[16'hFA00] = 8'hD8;
mem[16'hFA01] = 8'h62;
mem[16'hFA02] = 8'h5A;
mem[16'hFA03] = 8'h48;
mem[16'hFA04] = 8'h26;
mem[16'hFA05] = 8'h62;
mem[16'hFA06] = 8'h94;
mem[16'hFA07] = 8'h88;
mem[16'hFA08] = 8'h54;
mem[16'hFA09] = 8'h44;
mem[16'hFA0A] = 8'hC8;
mem[16'hFA0B] = 8'h54;
mem[16'hFA0C] = 8'h68;
mem[16'hFA0D] = 8'h44;
mem[16'hFA0E] = 8'hE8;
mem[16'hFA0F] = 8'h94;
mem[16'hFA10] = 8'h00;
mem[16'hFA11] = 8'hB4;
mem[16'hFA12] = 8'h08;
mem[16'hFA13] = 8'h84;
mem[16'hFA14] = 8'h74;
mem[16'hFA15] = 8'hB4;
mem[16'hFA16] = 8'h28;
mem[16'hFA17] = 8'h6E;
mem[16'hFA18] = 8'h74;
mem[16'hFA19] = 8'hF4;
mem[16'hFA1A] = 8'hCC;
mem[16'hFA1B] = 8'h4A;
mem[16'hFA1C] = 8'h72;
mem[16'hFA1D] = 8'hF2;
mem[16'hFA1E] = 8'hA4;
mem[16'hFA1F] = 8'h8A;
mem[16'hFA20] = 8'h00;
mem[16'hFA21] = 8'hAA;
mem[16'hFA22] = 8'hA2;
mem[16'hFA23] = 8'hA2;
mem[16'hFA24] = 8'h74;
mem[16'hFA25] = 8'h74;
mem[16'hFA26] = 8'h74;
mem[16'hFA27] = 8'h72;
mem[16'hFA28] = 8'h44;
mem[16'hFA29] = 8'h68;
mem[16'hFA2A] = 8'hB2;
mem[16'hFA2B] = 8'h32;
mem[16'hFA2C] = 8'hB2;
mem[16'hFA2D] = 8'h00;
mem[16'hFA2E] = 8'h22;
mem[16'hFA2F] = 8'h00;
mem[16'hFA30] = 8'h1A;
mem[16'hFA31] = 8'h1A;
mem[16'hFA32] = 8'h26;
mem[16'hFA33] = 8'h26;
mem[16'hFA34] = 8'h72;
mem[16'hFA35] = 8'h72;
mem[16'hFA36] = 8'h88;
mem[16'hFA37] = 8'hC8;
mem[16'hFA38] = 8'hC4;
mem[16'hFA39] = 8'hCA;
mem[16'hFA3A] = 8'h26;
mem[16'hFA3B] = 8'h48;
mem[16'hFA3C] = 8'h44;
mem[16'hFA3D] = 8'h44;
mem[16'hFA3E] = 8'hA2;
mem[16'hFA3F] = 8'hC8;
mem[16'hFA40] = 8'h85;
mem[16'hFA41] = 8'h45;
mem[16'hFA42] = 8'h68;
mem[16'hFA43] = 8'h48;
mem[16'hFA44] = 8'h0A;
mem[16'hFA45] = 8'h0A;
mem[16'hFA46] = 8'h0A;
mem[16'hFA47] = 8'h30;
mem[16'hFA48] = 8'h03;
mem[16'hFA49] = 8'h6C;
mem[16'hFA4A] = 8'hFE;
mem[16'hFA4B] = 8'h03;
mem[16'hFA4C] = 8'h28;
mem[16'hFA4D] = 8'h20;
mem[16'hFA4E] = 8'h4C;
mem[16'hFA4F] = 8'hFF;
mem[16'hFA50] = 8'h68;
mem[16'hFA51] = 8'h85;
mem[16'hFA52] = 8'h3A;
mem[16'hFA53] = 8'h68;
mem[16'hFA54] = 8'h85;
mem[16'hFA55] = 8'h3B;
mem[16'hFA56] = 8'h6C;
mem[16'hFA57] = 8'hF0;
mem[16'hFA58] = 8'h03;
mem[16'hFA59] = 8'h20;
mem[16'hFA5A] = 8'h82;
mem[16'hFA5B] = 8'hF8;
mem[16'hFA5C] = 8'h20;
mem[16'hFA5D] = 8'hDA;
mem[16'hFA5E] = 8'hFA;
mem[16'hFA5F] = 8'h4C;
mem[16'hFA60] = 8'h65;
mem[16'hFA61] = 8'hFF;
mem[16'hFA62] = 8'hD8;
mem[16'hFA63] = 8'h20;
mem[16'hFA64] = 8'h84;
mem[16'hFA65] = 8'hFE;
mem[16'hFA66] = 8'h20;
mem[16'hFA67] = 8'h2F;
mem[16'hFA68] = 8'hFB;
mem[16'hFA69] = 8'h20;
mem[16'hFA6A] = 8'h93;
mem[16'hFA6B] = 8'hFE;
mem[16'hFA6C] = 8'h20;
mem[16'hFA6D] = 8'h89;
mem[16'hFA6E] = 8'hFE;
mem[16'hFA6F] = 8'hAD;
mem[16'hFA70] = 8'h58;
mem[16'hFA71] = 8'hC0;
mem[16'hFA72] = 8'hAD;
mem[16'hFA73] = 8'h5A;
mem[16'hFA74] = 8'hC0;
mem[16'hFA75] = 8'hA0;
mem[16'hFA76] = 8'h05;
mem[16'hFA77] = 8'h20;
mem[16'hFA78] = 8'hB4;
mem[16'hFA79] = 8'hFB;
mem[16'hFA7A] = 8'hEA;
mem[16'hFA7B] = 8'hAD;
mem[16'hFA7C] = 8'hFF;
mem[16'hFA7D] = 8'hCF;
mem[16'hFA7E] = 8'h2C;
mem[16'hFA7F] = 8'h10;
mem[16'hFA80] = 8'hC0;
mem[16'hFA81] = 8'hD8;
mem[16'hFA82] = 8'h20;
mem[16'hFA83] = 8'h3A;
mem[16'hFA84] = 8'hFF;
mem[16'hFA85] = 8'hAD;
mem[16'hFA86] = 8'hF3;
mem[16'hFA87] = 8'h03;
mem[16'hFA88] = 8'h49;
mem[16'hFA89] = 8'hA5;
mem[16'hFA8A] = 8'hCD;
mem[16'hFA8B] = 8'hF4;
mem[16'hFA8C] = 8'h03;
mem[16'hFA8D] = 8'hD0;
mem[16'hFA8E] = 8'h17;
mem[16'hFA8F] = 8'hAD;
mem[16'hFA90] = 8'hF2;
mem[16'hFA91] = 8'h03;
mem[16'hFA92] = 8'hD0;
mem[16'hFA93] = 8'h0F;
mem[16'hFA94] = 8'hA9;
mem[16'hFA95] = 8'hE0;
mem[16'hFA96] = 8'hCD;
mem[16'hFA97] = 8'hF3;
mem[16'hFA98] = 8'h03;
mem[16'hFA99] = 8'hD0;
mem[16'hFA9A] = 8'h08;
mem[16'hFA9B] = 8'hA0;
mem[16'hFA9C] = 8'h03;
mem[16'hFA9D] = 8'h8C;
mem[16'hFA9E] = 8'hF2;
mem[16'hFA9F] = 8'h03;
mem[16'hFAA0] = 8'h4C;
mem[16'hFAA1] = 8'h00;
mem[16'hFAA2] = 8'hE0;
mem[16'hFAA3] = 8'h6C;
mem[16'hFAA4] = 8'hF2;
mem[16'hFAA5] = 8'h03;
mem[16'hFAA6] = 8'h20;
mem[16'hFAA7] = 8'h60;
mem[16'hFAA8] = 8'hFB;
mem[16'hFAA9] = 8'hA2;
mem[16'hFAAA] = 8'h05;
mem[16'hFAAB] = 8'hBD;
mem[16'hFAAC] = 8'hFC;
mem[16'hFAAD] = 8'hFA;
mem[16'hFAAE] = 8'h9D;
mem[16'hFAAF] = 8'hEF;
mem[16'hFAB0] = 8'h03;
mem[16'hFAB1] = 8'hCA;
mem[16'hFAB2] = 8'hD0;
mem[16'hFAB3] = 8'hF7;
mem[16'hFAB4] = 8'hA9;
mem[16'hFAB5] = 8'hC8;
mem[16'hFAB6] = 8'h86;
mem[16'hFAB7] = 8'h00;
mem[16'hFAB8] = 8'h85;
mem[16'hFAB9] = 8'h01;
mem[16'hFABA] = 8'hA0;
mem[16'hFABB] = 8'h07;
mem[16'hFABC] = 8'hC6;
mem[16'hFABD] = 8'h01;
mem[16'hFABE] = 8'hA5;
mem[16'hFABF] = 8'h01;
mem[16'hFAC0] = 8'hC9;
mem[16'hFAC1] = 8'hC0;
mem[16'hFAC2] = 8'hF0;
mem[16'hFAC3] = 8'hD7;
mem[16'hFAC4] = 8'h8D;
mem[16'hFAC5] = 8'hF8;
mem[16'hFAC6] = 8'h07;
mem[16'hFAC7] = 8'hB1;
mem[16'hFAC8] = 8'h00;
mem[16'hFAC9] = 8'hD9;
mem[16'hFACA] = 8'h01;
mem[16'hFACB] = 8'hFB;
mem[16'hFACC] = 8'hD0;
mem[16'hFACD] = 8'hEC;
mem[16'hFACE] = 8'h88;
mem[16'hFACF] = 8'h88;
mem[16'hFAD0] = 8'h10;
mem[16'hFAD1] = 8'hF5;
mem[16'hFAD2] = 8'h6C;
mem[16'hFAD3] = 8'h00;
mem[16'hFAD4] = 8'h00;
mem[16'hFAD5] = 8'hEA;
mem[16'hFAD6] = 8'hEA;
mem[16'hFAD7] = 8'h20;
mem[16'hFAD8] = 8'h8E;
mem[16'hFAD9] = 8'hFD;
mem[16'hFADA] = 8'hA9;
mem[16'hFADB] = 8'h45;
mem[16'hFADC] = 8'h85;
mem[16'hFADD] = 8'h40;
mem[16'hFADE] = 8'hA9;
mem[16'hFADF] = 8'h00;
mem[16'hFAE0] = 8'h85;
mem[16'hFAE1] = 8'h41;
mem[16'hFAE2] = 8'hA2;
mem[16'hFAE3] = 8'hFB;
mem[16'hFAE4] = 8'hA9;
mem[16'hFAE5] = 8'hA0;
mem[16'hFAE6] = 8'h20;
mem[16'hFAE7] = 8'hED;
mem[16'hFAE8] = 8'hFD;
mem[16'hFAE9] = 8'hBD;
mem[16'hFAEA] = 8'h1E;
mem[16'hFAEB] = 8'hFA;
mem[16'hFAEC] = 8'h20;
mem[16'hFAED] = 8'hED;
mem[16'hFAEE] = 8'hFD;
mem[16'hFAEF] = 8'hA9;
mem[16'hFAF0] = 8'hBD;
mem[16'hFAF1] = 8'h20;
mem[16'hFAF2] = 8'hED;
mem[16'hFAF3] = 8'hFD;
mem[16'hFAF4] = 8'hB5;
mem[16'hFAF5] = 8'h4A;
mem[16'hFAF6] = 8'h20;
mem[16'hFAF7] = 8'hDA;
mem[16'hFAF8] = 8'hFD;
mem[16'hFAF9] = 8'hE8;
mem[16'hFAFA] = 8'h30;
mem[16'hFAFB] = 8'hE8;
mem[16'hFAFC] = 8'h60;
mem[16'hFAFD] = 8'h59;
mem[16'hFAFE] = 8'hFA;
mem[16'hFAFF] = 8'h00;
mem[16'hFB00] = 8'hE0;
mem[16'hFB01] = 8'h45;
mem[16'hFB02] = 8'h20;
mem[16'hFB03] = 8'hFF;
mem[16'hFB04] = 8'h00;
mem[16'hFB05] = 8'hFF;
mem[16'hFB06] = 8'h03;
mem[16'hFB07] = 8'hFF;
mem[16'hFB08] = 8'h3C;
mem[16'hFB09] = 8'hC1;
mem[16'hFB0A] = 8'hF0;
mem[16'hFB0B] = 8'hF0;
mem[16'hFB0C] = 8'hEC;
mem[16'hFB0D] = 8'hE5;
mem[16'hFB0E] = 8'hA0;
mem[16'hFB0F] = 8'hDD;
mem[16'hFB10] = 8'hDB;
mem[16'hFB11] = 8'hC4;
mem[16'hFB12] = 8'hC2;
mem[16'hFB13] = 8'hC1;
mem[16'hFB14] = 8'hFF;
mem[16'hFB15] = 8'hC3;
mem[16'hFB16] = 8'hFF;
mem[16'hFB17] = 8'hFF;
mem[16'hFB18] = 8'hFF;
mem[16'hFB19] = 8'hC1;
mem[16'hFB1A] = 8'hD8;
mem[16'hFB1B] = 8'hD9;
mem[16'hFB1C] = 8'hD0;
mem[16'hFB1D] = 8'hD3;
mem[16'hFB1E] = 8'hAD;
mem[16'hFB1F] = 8'h70;
mem[16'hFB20] = 8'hC0;
mem[16'hFB21] = 8'hA0;
mem[16'hFB22] = 8'h00;
mem[16'hFB23] = 8'hEA;
mem[16'hFB24] = 8'hEA;
mem[16'hFB25] = 8'hBD;
mem[16'hFB26] = 8'h64;
mem[16'hFB27] = 8'hC0;
mem[16'hFB28] = 8'h10;
mem[16'hFB29] = 8'h04;
mem[16'hFB2A] = 8'hC8;
mem[16'hFB2B] = 8'hD0;
mem[16'hFB2C] = 8'hF8;
mem[16'hFB2D] = 8'h88;
mem[16'hFB2E] = 8'h60;
mem[16'hFB2F] = 8'hA9;
mem[16'hFB30] = 8'h00;
mem[16'hFB31] = 8'h85;
mem[16'hFB32] = 8'h48;
mem[16'hFB33] = 8'hAD;
mem[16'hFB34] = 8'h56;
mem[16'hFB35] = 8'hC0;
mem[16'hFB36] = 8'hAD;
mem[16'hFB37] = 8'h54;
mem[16'hFB38] = 8'hC0;
mem[16'hFB39] = 8'hAD;
mem[16'hFB3A] = 8'h51;
mem[16'hFB3B] = 8'hC0;
mem[16'hFB3C] = 8'hA9;
mem[16'hFB3D] = 8'h00;
mem[16'hFB3E] = 8'hF0;
mem[16'hFB3F] = 8'h0B;
mem[16'hFB40] = 8'hAD;
mem[16'hFB41] = 8'h50;
mem[16'hFB42] = 8'hC0;
mem[16'hFB43] = 8'hAD;
mem[16'hFB44] = 8'h53;
mem[16'hFB45] = 8'hC0;
mem[16'hFB46] = 8'h20;
mem[16'hFB47] = 8'h36;
mem[16'hFB48] = 8'hF8;
mem[16'hFB49] = 8'hA9;
mem[16'hFB4A] = 8'h14;
mem[16'hFB4B] = 8'h85;
mem[16'hFB4C] = 8'h22;
mem[16'hFB4D] = 8'hA9;
mem[16'hFB4E] = 8'h00;
mem[16'hFB4F] = 8'h85;
mem[16'hFB50] = 8'h20;
mem[16'hFB51] = 8'hA0;
mem[16'hFB52] = 8'h08;
mem[16'hFB53] = 8'hD0;
mem[16'hFB54] = 8'h5F;
mem[16'hFB55] = 8'hA9;
mem[16'hFB56] = 8'h18;
mem[16'hFB57] = 8'h85;
mem[16'hFB58] = 8'h23;
mem[16'hFB59] = 8'hA9;
mem[16'hFB5A] = 8'h17;
mem[16'hFB5B] = 8'h85;
mem[16'hFB5C] = 8'h25;
mem[16'hFB5D] = 8'h4C;
mem[16'hFB5E] = 8'h22;
mem[16'hFB5F] = 8'hFC;
mem[16'hFB60] = 8'h20;
mem[16'hFB61] = 8'h58;
mem[16'hFB62] = 8'hFC;
mem[16'hFB63] = 8'hA0;
mem[16'hFB64] = 8'h08;
mem[16'hFB65] = 8'hB9;
mem[16'hFB66] = 8'h08;
mem[16'hFB67] = 8'hFB;
mem[16'hFB68] = 8'h99;
mem[16'hFB69] = 8'h0E;
mem[16'hFB6A] = 8'h04;
mem[16'hFB6B] = 8'h88;
mem[16'hFB6C] = 8'hD0;
mem[16'hFB6D] = 8'hF7;
mem[16'hFB6E] = 8'h60;
mem[16'hFB6F] = 8'hAD;
mem[16'hFB70] = 8'hF3;
mem[16'hFB71] = 8'h03;
mem[16'hFB72] = 8'h49;
mem[16'hFB73] = 8'hA5;
mem[16'hFB74] = 8'h8D;
mem[16'hFB75] = 8'hF4;
mem[16'hFB76] = 8'h03;
mem[16'hFB77] = 8'h60;
mem[16'hFB78] = 8'hC9;
mem[16'hFB79] = 8'h8D;
mem[16'hFB7A] = 8'hD0;
mem[16'hFB7B] = 8'h18;
mem[16'hFB7C] = 8'hAC;
mem[16'hFB7D] = 8'h00;
mem[16'hFB7E] = 8'hC0;
mem[16'hFB7F] = 8'h10;
mem[16'hFB80] = 8'h13;
mem[16'hFB81] = 8'hC0;
mem[16'hFB82] = 8'h93;
mem[16'hFB83] = 8'hD0;
mem[16'hFB84] = 8'h0F;
mem[16'hFB85] = 8'h2C;
mem[16'hFB86] = 8'h10;
mem[16'hFB87] = 8'hC0;
mem[16'hFB88] = 8'hAC;
mem[16'hFB89] = 8'h00;
mem[16'hFB8A] = 8'hC0;
mem[16'hFB8B] = 8'h10;
mem[16'hFB8C] = 8'hFB;
mem[16'hFB8D] = 8'hC0;
mem[16'hFB8E] = 8'h83;
mem[16'hFB8F] = 8'hF0;
mem[16'hFB90] = 8'h03;
mem[16'hFB91] = 8'h2C;
mem[16'hFB92] = 8'h10;
mem[16'hFB93] = 8'hC0;
mem[16'hFB94] = 8'h4C;
mem[16'hFB95] = 8'hFD;
mem[16'hFB96] = 8'hFB;
mem[16'hFB97] = 8'h38;
mem[16'hFB98] = 8'h4C;
mem[16'hFB99] = 8'h2C;
mem[16'hFB9A] = 8'hFC;
mem[16'hFB9B] = 8'hA8;
mem[16'hFB9C] = 8'hB9;
mem[16'hFB9D] = 8'h48;
mem[16'hFB9E] = 8'hFA;
mem[16'hFB9F] = 8'h20;
mem[16'hFBA0] = 8'h97;
mem[16'hFBA1] = 8'hFB;
mem[16'hFBA2] = 8'h20;
mem[16'hFBA3] = 8'h21;
mem[16'hFBA4] = 8'hFD;
mem[16'hFBA5] = 8'hC9;
mem[16'hFBA6] = 8'hCE;
mem[16'hFBA7] = 8'hB0;
mem[16'hFBA8] = 8'hEE;
mem[16'hFBA9] = 8'hC9;
mem[16'hFBAA] = 8'hC9;
mem[16'hFBAB] = 8'h90;
mem[16'hFBAC] = 8'hEA;
mem[16'hFBAD] = 8'hC9;
mem[16'hFBAE] = 8'hCC;
mem[16'hFBAF] = 8'hF0;
mem[16'hFBB0] = 8'hE6;
mem[16'hFBB1] = 8'hD0;
mem[16'hFBB2] = 8'hE8;
mem[16'hFBB3] = 8'h06;
mem[16'hFBB4] = 8'h08;
mem[16'hFBB5] = 8'h78;
mem[16'hFBB6] = 8'h2C;
mem[16'hFBB7] = 8'h15;
mem[16'hFBB8] = 8'hC0;
mem[16'hFBB9] = 8'h08;
mem[16'hFBBA] = 8'h8D;
mem[16'hFBBB] = 8'h07;
mem[16'hFBBC] = 8'hC0;
mem[16'hFBBD] = 8'h4C;
mem[16'hFBBE] = 8'h00;
mem[16'hFBBF] = 8'hC1;
mem[16'hFBC0] = 8'hEA;
mem[16'hFBC1] = 8'h48;
mem[16'hFBC2] = 8'h4A;
mem[16'hFBC3] = 8'h29;
mem[16'hFBC4] = 8'h03;
mem[16'hFBC5] = 8'h09;
mem[16'hFBC6] = 8'h04;
mem[16'hFBC7] = 8'h85;
mem[16'hFBC8] = 8'h29;
mem[16'hFBC9] = 8'h68;
mem[16'hFBCA] = 8'h29;
mem[16'hFBCB] = 8'h18;
mem[16'hFBCC] = 8'h90;
mem[16'hFBCD] = 8'h02;
mem[16'hFBCE] = 8'h69;
mem[16'hFBCF] = 8'h7F;
mem[16'hFBD0] = 8'h85;
mem[16'hFBD1] = 8'h28;
mem[16'hFBD2] = 8'h0A;
mem[16'hFBD3] = 8'h0A;
mem[16'hFBD4] = 8'h05;
mem[16'hFBD5] = 8'h28;
mem[16'hFBD6] = 8'h85;
mem[16'hFBD7] = 8'h28;
mem[16'hFBD8] = 8'h60;
mem[16'hFBD9] = 8'hC9;
mem[16'hFBDA] = 8'h87;
mem[16'hFBDB] = 8'hD0;
mem[16'hFBDC] = 8'h12;
mem[16'hFBDD] = 8'hA9;
mem[16'hFBDE] = 8'h40;
mem[16'hFBDF] = 8'h20;
mem[16'hFBE0] = 8'hA8;
mem[16'hFBE1] = 8'hFC;
mem[16'hFBE2] = 8'hA0;
mem[16'hFBE3] = 8'hC0;
mem[16'hFBE4] = 8'hA9;
mem[16'hFBE5] = 8'h0C;
mem[16'hFBE6] = 8'h20;
mem[16'hFBE7] = 8'hA8;
mem[16'hFBE8] = 8'hFC;
mem[16'hFBE9] = 8'hAD;
mem[16'hFBEA] = 8'h30;
mem[16'hFBEB] = 8'hC0;
mem[16'hFBEC] = 8'h88;
mem[16'hFBED] = 8'hD0;
mem[16'hFBEE] = 8'hF5;
mem[16'hFBEF] = 8'h60;
mem[16'hFBF0] = 8'hA4;
mem[16'hFBF1] = 8'h24;
mem[16'hFBF2] = 8'h91;
mem[16'hFBF3] = 8'h28;
mem[16'hFBF4] = 8'hE6;
mem[16'hFBF5] = 8'h24;
mem[16'hFBF6] = 8'hA5;
mem[16'hFBF7] = 8'h24;
mem[16'hFBF8] = 8'hC5;
mem[16'hFBF9] = 8'h21;
mem[16'hFBFA] = 8'hB0;
mem[16'hFBFB] = 8'h66;
mem[16'hFBFC] = 8'h60;
mem[16'hFBFD] = 8'hC9;
mem[16'hFBFE] = 8'hA0;
mem[16'hFBFF] = 8'hB0;
mem[16'hFC00] = 8'hEF;
mem[16'hFC01] = 8'hA8;
mem[16'hFC02] = 8'h10;
mem[16'hFC03] = 8'hEC;
mem[16'hFC04] = 8'hC9;
mem[16'hFC05] = 8'h8D;
mem[16'hFC06] = 8'hF0;
mem[16'hFC07] = 8'h5A;
mem[16'hFC08] = 8'hC9;
mem[16'hFC09] = 8'h8A;
mem[16'hFC0A] = 8'hF0;
mem[16'hFC0B] = 8'h5A;
mem[16'hFC0C] = 8'hC9;
mem[16'hFC0D] = 8'h88;
mem[16'hFC0E] = 8'hD0;
mem[16'hFC0F] = 8'hC9;
mem[16'hFC10] = 8'hC6;
mem[16'hFC11] = 8'h24;
mem[16'hFC12] = 8'h10;
mem[16'hFC13] = 8'hE8;
mem[16'hFC14] = 8'hA5;
mem[16'hFC15] = 8'h21;
mem[16'hFC16] = 8'h85;
mem[16'hFC17] = 8'h24;
mem[16'hFC18] = 8'hC6;
mem[16'hFC19] = 8'h24;
mem[16'hFC1A] = 8'hA5;
mem[16'hFC1B] = 8'h22;
mem[16'hFC1C] = 8'hC5;
mem[16'hFC1D] = 8'h25;
mem[16'hFC1E] = 8'hB0;
mem[16'hFC1F] = 8'h0B;
mem[16'hFC20] = 8'hC6;
mem[16'hFC21] = 8'h25;
mem[16'hFC22] = 8'hA5;
mem[16'hFC23] = 8'h25;
mem[16'hFC24] = 8'h20;
mem[16'hFC25] = 8'hC1;
mem[16'hFC26] = 8'hFB;
mem[16'hFC27] = 8'h65;
mem[16'hFC28] = 8'h20;
mem[16'hFC29] = 8'h85;
mem[16'hFC2A] = 8'h28;
mem[16'hFC2B] = 8'h60;
mem[16'hFC2C] = 8'h49;
mem[16'hFC2D] = 8'hC0;
mem[16'hFC2E] = 8'hF0;
mem[16'hFC2F] = 8'h28;
mem[16'hFC30] = 8'h69;
mem[16'hFC31] = 8'hFD;
mem[16'hFC32] = 8'h90;
mem[16'hFC33] = 8'hC0;
mem[16'hFC34] = 8'hF0;
mem[16'hFC35] = 8'hDA;
mem[16'hFC36] = 8'h69;
mem[16'hFC37] = 8'hFD;
mem[16'hFC38] = 8'h90;
mem[16'hFC39] = 8'h2C;
mem[16'hFC3A] = 8'hF0;
mem[16'hFC3B] = 8'hDE;
mem[16'hFC3C] = 8'h69;
mem[16'hFC3D] = 8'hFD;
mem[16'hFC3E] = 8'h90;
mem[16'hFC3F] = 8'h5C;
mem[16'hFC40] = 8'hD0;
mem[16'hFC41] = 8'hE9;
mem[16'hFC42] = 8'hA0;
mem[16'hFC43] = 8'h00;
mem[16'hFC44] = 8'hF0;
mem[16'hFC45] = 8'h2C;
mem[16'hFC46] = 8'hA8;
mem[16'hFC47] = 8'hC3;
mem[16'hFC48] = 8'hA9;
mem[16'hFC49] = 8'hA0;
mem[16'hFC4A] = 8'hB1;
mem[16'hFC4B] = 8'hB9;
mem[16'hFC4C] = 8'hB8;
mem[16'hFC4D] = 8'hB1;
mem[16'hFC4E] = 8'hAD;
mem[16'hFC4F] = 8'hB8;
mem[16'hFC50] = 8'hB2;
mem[16'hFC51] = 8'hAC;
mem[16'hFC52] = 8'hA0;
mem[16'hFC53] = 8'hC1;
mem[16'hFC54] = 8'hD0;
mem[16'hFC55] = 8'hD0;
mem[16'hFC56] = 8'hCC;
mem[16'hFC57] = 8'hC5;
mem[16'hFC58] = 8'hA0;
mem[16'hFC59] = 8'h01;
mem[16'hFC5A] = 8'hD0;
mem[16'hFC5B] = 8'h16;
mem[16'hFC5C] = 8'hD2;
mem[16'hFC5D] = 8'hC9;
mem[16'hFC5E] = 8'hC3;
mem[16'hFC5F] = 8'hCB;
mem[16'hFC60] = 8'hA0;
mem[16'hFC61] = 8'hC1;
mem[16'hFC62] = 8'hA9;
mem[16'hFC63] = 8'h00;
mem[16'hFC64] = 8'h85;
mem[16'hFC65] = 8'h24;
mem[16'hFC66] = 8'hE6;
mem[16'hFC67] = 8'h25;
mem[16'hFC68] = 8'hA5;
mem[16'hFC69] = 8'h25;
mem[16'hFC6A] = 8'hC5;
mem[16'hFC6B] = 8'h23;
mem[16'hFC6C] = 8'h90;
mem[16'hFC6D] = 8'hB6;
mem[16'hFC6E] = 8'hC6;
mem[16'hFC6F] = 8'h25;
mem[16'hFC70] = 8'hA0;
mem[16'hFC71] = 8'h02;
mem[16'hFC72] = 8'h4C;
mem[16'hFC73] = 8'hB4;
mem[16'hFC74] = 8'hFB;
mem[16'hFC75] = 8'h48;
mem[16'hFC76] = 8'hAD;
mem[16'hFC77] = 8'h18;
mem[16'hFC78] = 8'hC0;
mem[16'hFC79] = 8'h0A;
mem[16'hFC7A] = 8'h68;
mem[16'hFC7B] = 8'h2C;
mem[16'hFC7C] = 8'h1C;
mem[16'hFC7D] = 8'hC0;
mem[16'hFC7E] = 8'h08;
mem[16'hFC7F] = 8'h90;
mem[16'hFC80] = 8'h03;
mem[16'hFC81] = 8'h8D;
mem[16'hFC82] = 8'h54;
mem[16'hFC83] = 8'hC0;
mem[16'hFC84] = 8'h2C;
mem[16'hFC85] = 8'h15;
mem[16'hFC86] = 8'hC0;
mem[16'hFC87] = 8'h8D;
mem[16'hFC88] = 8'h06;
mem[16'hFC89] = 8'hC0;
mem[16'hFC8A] = 8'h58;
mem[16'hFC8B] = 8'h78;
mem[16'hFC8C] = 8'h10;
mem[16'hFC8D] = 8'h03;
mem[16'hFC8E] = 8'h8D;
mem[16'hFC8F] = 8'h07;
mem[16'hFC90] = 8'hC0;
mem[16'hFC91] = 8'h28;
mem[16'hFC92] = 8'h90;
mem[16'hFC93] = 8'h05;
mem[16'hFC94] = 8'h10;
mem[16'hFC95] = 8'h03;
mem[16'hFC96] = 8'h2C;
mem[16'hFC97] = 8'h55;
mem[16'hFC98] = 8'hC0;
mem[16'hFC99] = 8'h60;
mem[16'hFC9A] = 8'hEA;
mem[16'hFC9B] = 8'hEA;
mem[16'hFC9C] = 8'h18;
mem[16'hFC9D] = 8'hB0;
mem[16'hFC9E] = 8'h38;
mem[16'hFC9F] = 8'h84;
mem[16'hFCA0] = 8'h1F;
mem[16'hFCA1] = 8'hA0;
mem[16'hFCA2] = 8'h03;
mem[16'hFCA3] = 8'h90;
mem[16'hFCA4] = 8'hCD;
mem[16'hFCA5] = 8'hC8;
mem[16'hFCA6] = 8'hD0;
mem[16'hFCA7] = 8'hCA;
mem[16'hFCA8] = 8'h38;
mem[16'hFCA9] = 8'h48;
mem[16'hFCAA] = 8'hE9;
mem[16'hFCAB] = 8'h01;
mem[16'hFCAC] = 8'hD0;
mem[16'hFCAD] = 8'hFC;
mem[16'hFCAE] = 8'h68;
mem[16'hFCAF] = 8'hE9;
mem[16'hFCB0] = 8'h01;
mem[16'hFCB1] = 8'hD0;
mem[16'hFCB2] = 8'hF6;
mem[16'hFCB3] = 8'h60;
mem[16'hFCB4] = 8'hE6;
mem[16'hFCB5] = 8'h42;
mem[16'hFCB6] = 8'hD0;
mem[16'hFCB7] = 8'h02;
mem[16'hFCB8] = 8'hE6;
mem[16'hFCB9] = 8'h43;
mem[16'hFCBA] = 8'hA5;
mem[16'hFCBB] = 8'h3C;
mem[16'hFCBC] = 8'hC5;
mem[16'hFCBD] = 8'h3E;
mem[16'hFCBE] = 8'hA5;
mem[16'hFCBF] = 8'h3D;
mem[16'hFCC0] = 8'hE5;
mem[16'hFCC1] = 8'h3F;
mem[16'hFCC2] = 8'hE6;
mem[16'hFCC3] = 8'h3C;
mem[16'hFCC4] = 8'hD0;
mem[16'hFCC5] = 8'h02;
mem[16'hFCC6] = 8'hE6;
mem[16'hFCC7] = 8'h3D;
mem[16'hFCC8] = 8'h60;
mem[16'hFCC9] = 8'hA0;
mem[16'hFCCA] = 8'h4B;
mem[16'hFCCB] = 8'h20;
mem[16'hFCCC] = 8'hDB;
mem[16'hFCCD] = 8'hFC;
mem[16'hFCCE] = 8'hD0;
mem[16'hFCCF] = 8'hF9;
mem[16'hFCD0] = 8'h69;
mem[16'hFCD1] = 8'hFE;
mem[16'hFCD2] = 8'hB0;
mem[16'hFCD3] = 8'hF5;
mem[16'hFCD4] = 8'hA0;
mem[16'hFCD5] = 8'h21;
mem[16'hFCD6] = 8'h20;
mem[16'hFCD7] = 8'hDB;
mem[16'hFCD8] = 8'hFC;
mem[16'hFCD9] = 8'hC8;
mem[16'hFCDA] = 8'hC8;
mem[16'hFCDB] = 8'h88;
mem[16'hFCDC] = 8'hD0;
mem[16'hFCDD] = 8'hFD;
mem[16'hFCDE] = 8'h90;
mem[16'hFCDF] = 8'h05;
mem[16'hFCE0] = 8'hA0;
mem[16'hFCE1] = 8'h32;
mem[16'hFCE2] = 8'h88;
mem[16'hFCE3] = 8'hD0;
mem[16'hFCE4] = 8'hFD;
mem[16'hFCE5] = 8'hAC;
mem[16'hFCE6] = 8'h20;
mem[16'hFCE7] = 8'hC0;
mem[16'hFCE8] = 8'hA0;
mem[16'hFCE9] = 8'h2C;
mem[16'hFCEA] = 8'hCA;
mem[16'hFCEB] = 8'h60;
mem[16'hFCEC] = 8'hA2;
mem[16'hFCED] = 8'h08;
mem[16'hFCEE] = 8'h48;
mem[16'hFCEF] = 8'h20;
mem[16'hFCF0] = 8'hFA;
mem[16'hFCF1] = 8'hFC;
mem[16'hFCF2] = 8'h68;
mem[16'hFCF3] = 8'h2A;
mem[16'hFCF4] = 8'hA0;
mem[16'hFCF5] = 8'h3A;
mem[16'hFCF6] = 8'hCA;
mem[16'hFCF7] = 8'hD0;
mem[16'hFCF8] = 8'hF5;
mem[16'hFCF9] = 8'h60;
mem[16'hFCFA] = 8'h20;
mem[16'hFCFB] = 8'hFD;
mem[16'hFCFC] = 8'hFC;
mem[16'hFCFD] = 8'h88;
mem[16'hFCFE] = 8'hAD;
mem[16'hFCFF] = 8'h60;
mem[16'hFD00] = 8'hC0;
mem[16'hFD01] = 8'h45;
mem[16'hFD02] = 8'h2F;
mem[16'hFD03] = 8'h10;
mem[16'hFD04] = 8'hF8;
mem[16'hFD05] = 8'h45;
mem[16'hFD06] = 8'h2F;
mem[16'hFD07] = 8'h85;
mem[16'hFD08] = 8'h2F;
mem[16'hFD09] = 8'hC0;
mem[16'hFD0A] = 8'h80;
mem[16'hFD0B] = 8'h60;
mem[16'hFD0C] = 8'hA4;
mem[16'hFD0D] = 8'h24;
mem[16'hFD0E] = 8'hB1;
mem[16'hFD0F] = 8'h28;
mem[16'hFD10] = 8'h48;
mem[16'hFD11] = 8'h29;
mem[16'hFD12] = 8'h3F;
mem[16'hFD13] = 8'h09;
mem[16'hFD14] = 8'h40;
mem[16'hFD15] = 8'h91;
mem[16'hFD16] = 8'h28;
mem[16'hFD17] = 8'h68;
mem[16'hFD18] = 8'h6C;
mem[16'hFD19] = 8'h38;
mem[16'hFD1A] = 8'h00;
mem[16'hFD1B] = 8'hA0;
mem[16'hFD1C] = 8'h06;
mem[16'hFD1D] = 8'h4C;
mem[16'hFD1E] = 8'hB4;
mem[16'hFD1F] = 8'hFB;
mem[16'hFD20] = 8'hEA;
mem[16'hFD21] = 8'h20;
mem[16'hFD22] = 8'h0C;
mem[16'hFD23] = 8'hFD;
mem[16'hFD24] = 8'hA0;
mem[16'hFD25] = 8'h07;
mem[16'hFD26] = 8'h4C;
mem[16'hFD27] = 8'hB4;
mem[16'hFD28] = 8'hFB;
mem[16'hFD29] = 8'h8D;
mem[16'hFD2A] = 8'h06;
mem[16'hFD2B] = 8'hC0;
mem[16'hFD2C] = 8'h28;
mem[16'hFD2D] = 8'h60;
mem[16'hFD2E] = 8'h60;
mem[16'hFD2F] = 8'h20;
mem[16'hFD30] = 8'h21;
mem[16'hFD31] = 8'hFD;
mem[16'hFD32] = 8'h20;
mem[16'hFD33] = 8'hA5;
mem[16'hFD34] = 8'hFB;
mem[16'hFD35] = 8'h20;
mem[16'hFD36] = 8'h0C;
mem[16'hFD37] = 8'hFD;
mem[16'hFD38] = 8'hC9;
mem[16'hFD39] = 8'h9B;
mem[16'hFD3A] = 8'hF0;
mem[16'hFD3B] = 8'hF3;
mem[16'hFD3C] = 8'h60;
mem[16'hFD3D] = 8'hA5;
mem[16'hFD3E] = 8'h32;
mem[16'hFD3F] = 8'h48;
mem[16'hFD40] = 8'hA9;
mem[16'hFD41] = 8'hFF;
mem[16'hFD42] = 8'hEA;
mem[16'hFD43] = 8'hEA;
mem[16'hFD44] = 8'hBD;
mem[16'hFD45] = 8'h00;
mem[16'hFD46] = 8'h02;
mem[16'hFD47] = 8'h20;
mem[16'hFD48] = 8'hED;
mem[16'hFD49] = 8'hFD;
mem[16'hFD4A] = 8'h68;
mem[16'hFD4B] = 8'h85;
mem[16'hFD4C] = 8'h32;
mem[16'hFD4D] = 8'hBD;
mem[16'hFD4E] = 8'h00;
mem[16'hFD4F] = 8'h02;
mem[16'hFD50] = 8'hC9;
mem[16'hFD51] = 8'h88;
mem[16'hFD52] = 8'hF0;
mem[16'hFD53] = 8'h1D;
mem[16'hFD54] = 8'hC9;
mem[16'hFD55] = 8'h98;
mem[16'hFD56] = 8'hF0;
mem[16'hFD57] = 8'h0A;
mem[16'hFD58] = 8'hE0;
mem[16'hFD59] = 8'hF8;
mem[16'hFD5A] = 8'h90;
mem[16'hFD5B] = 8'h03;
mem[16'hFD5C] = 8'h20;
mem[16'hFD5D] = 8'h3A;
mem[16'hFD5E] = 8'hFF;
mem[16'hFD5F] = 8'hE8;
mem[16'hFD60] = 8'hD0;
mem[16'hFD61] = 8'h13;
mem[16'hFD62] = 8'hA9;
mem[16'hFD63] = 8'hDC;
mem[16'hFD64] = 8'h20;
mem[16'hFD65] = 8'hED;
mem[16'hFD66] = 8'hFD;
mem[16'hFD67] = 8'h20;
mem[16'hFD68] = 8'h8E;
mem[16'hFD69] = 8'hFD;
mem[16'hFD6A] = 8'hA5;
mem[16'hFD6B] = 8'h33;
mem[16'hFD6C] = 8'h20;
mem[16'hFD6D] = 8'hED;
mem[16'hFD6E] = 8'hFD;
mem[16'hFD6F] = 8'hA2;
mem[16'hFD70] = 8'h01;
mem[16'hFD71] = 8'h8A;
mem[16'hFD72] = 8'hF0;
mem[16'hFD73] = 8'hF3;
mem[16'hFD74] = 8'hCA;
mem[16'hFD75] = 8'h20;
mem[16'hFD76] = 8'h35;
mem[16'hFD77] = 8'hFD;
mem[16'hFD78] = 8'hC9;
mem[16'hFD79] = 8'h95;
mem[16'hFD7A] = 8'hD0;
mem[16'hFD7B] = 8'h02;
mem[16'hFD7C] = 8'hB1;
mem[16'hFD7D] = 8'h28;
mem[16'hFD7E] = 8'hC9;
mem[16'hFD7F] = 8'hE0;
mem[16'hFD80] = 8'h90;
mem[16'hFD81] = 8'h02;
mem[16'hFD82] = 8'h29;
mem[16'hFD83] = 8'hFF;
mem[16'hFD84] = 8'h9D;
mem[16'hFD85] = 8'h00;
mem[16'hFD86] = 8'h02;
mem[16'hFD87] = 8'hC9;
mem[16'hFD88] = 8'h8D;
mem[16'hFD89] = 8'hD0;
mem[16'hFD8A] = 8'hB2;
mem[16'hFD8B] = 8'h20;
mem[16'hFD8C] = 8'h9C;
mem[16'hFD8D] = 8'hFC;
mem[16'hFD8E] = 8'hA9;
mem[16'hFD8F] = 8'h8D;
mem[16'hFD90] = 8'hD0;
mem[16'hFD91] = 8'h5B;
mem[16'hFD92] = 8'hA4;
mem[16'hFD93] = 8'h3D;
mem[16'hFD94] = 8'hA6;
mem[16'hFD95] = 8'h3C;
mem[16'hFD96] = 8'h20;
mem[16'hFD97] = 8'h8E;
mem[16'hFD98] = 8'hFD;
mem[16'hFD99] = 8'h20;
mem[16'hFD9A] = 8'h40;
mem[16'hFD9B] = 8'hF9;
mem[16'hFD9C] = 8'hA0;
mem[16'hFD9D] = 8'h00;
mem[16'hFD9E] = 8'hA9;
mem[16'hFD9F] = 8'hAD;
mem[16'hFDA0] = 8'h4C;
mem[16'hFDA1] = 8'hED;
mem[16'hFDA2] = 8'hFD;
mem[16'hFDA3] = 8'hA5;
mem[16'hFDA4] = 8'h3C;
mem[16'hFDA5] = 8'h09;
mem[16'hFDA6] = 8'h07;
mem[16'hFDA7] = 8'h85;
mem[16'hFDA8] = 8'h3E;
mem[16'hFDA9] = 8'hA5;
mem[16'hFDAA] = 8'h3D;
mem[16'hFDAB] = 8'h85;
mem[16'hFDAC] = 8'h3F;
mem[16'hFDAD] = 8'hA5;
mem[16'hFDAE] = 8'h3C;
mem[16'hFDAF] = 8'h29;
mem[16'hFDB0] = 8'h07;
mem[16'hFDB1] = 8'hD0;
mem[16'hFDB2] = 8'h03;
mem[16'hFDB3] = 8'h20;
mem[16'hFDB4] = 8'h92;
mem[16'hFDB5] = 8'hFD;
mem[16'hFDB6] = 8'hA9;
mem[16'hFDB7] = 8'hA0;
mem[16'hFDB8] = 8'h20;
mem[16'hFDB9] = 8'hED;
mem[16'hFDBA] = 8'hFD;
mem[16'hFDBB] = 8'hB1;
mem[16'hFDBC] = 8'h3C;
mem[16'hFDBD] = 8'h20;
mem[16'hFDBE] = 8'hDA;
mem[16'hFDBF] = 8'hFD;
mem[16'hFDC0] = 8'h20;
mem[16'hFDC1] = 8'hBA;
mem[16'hFDC2] = 8'hFC;
mem[16'hFDC3] = 8'h90;
mem[16'hFDC4] = 8'hE8;
mem[16'hFDC5] = 8'h60;
mem[16'hFDC6] = 8'h4A;
mem[16'hFDC7] = 8'h90;
mem[16'hFDC8] = 8'hEA;
mem[16'hFDC9] = 8'h4A;
mem[16'hFDCA] = 8'h4A;
mem[16'hFDCB] = 8'hA5;
mem[16'hFDCC] = 8'h3E;
mem[16'hFDCD] = 8'h90;
mem[16'hFDCE] = 8'h02;
mem[16'hFDCF] = 8'h49;
mem[16'hFDD0] = 8'hFF;
mem[16'hFDD1] = 8'h65;
mem[16'hFDD2] = 8'h3C;
mem[16'hFDD3] = 8'h48;
mem[16'hFDD4] = 8'hA9;
mem[16'hFDD5] = 8'hBD;
mem[16'hFDD6] = 8'h20;
mem[16'hFDD7] = 8'hED;
mem[16'hFDD8] = 8'hFD;
mem[16'hFDD9] = 8'h68;
mem[16'hFDDA] = 8'h48;
mem[16'hFDDB] = 8'h4A;
mem[16'hFDDC] = 8'h4A;
mem[16'hFDDD] = 8'h4A;
mem[16'hFDDE] = 8'h4A;
mem[16'hFDDF] = 8'h20;
mem[16'hFDE0] = 8'hE5;
mem[16'hFDE1] = 8'hFD;
mem[16'hFDE2] = 8'h68;
mem[16'hFDE3] = 8'h29;
mem[16'hFDE4] = 8'h0F;
mem[16'hFDE5] = 8'h09;
mem[16'hFDE6] = 8'hB0;
mem[16'hFDE7] = 8'hC9;
mem[16'hFDE8] = 8'hBA;
mem[16'hFDE9] = 8'h90;
mem[16'hFDEA] = 8'h02;
mem[16'hFDEB] = 8'h69;
mem[16'hFDEC] = 8'h06;
mem[16'hFDED] = 8'h6C;
mem[16'hFDEE] = 8'h36;
mem[16'hFDEF] = 8'h00;
mem[16'hFDF0] = 8'hC9;
mem[16'hFDF1] = 8'hA0;
mem[16'hFDF2] = 8'h90;
mem[16'hFDF3] = 8'h02;
mem[16'hFDF4] = 8'h25;
mem[16'hFDF5] = 8'h32;
mem[16'hFDF6] = 8'h84;
mem[16'hFDF7] = 8'h35;
mem[16'hFDF8] = 8'h48;
mem[16'hFDF9] = 8'h20;
mem[16'hFDFA] = 8'h78;
mem[16'hFDFB] = 8'hFB;
mem[16'hFDFC] = 8'h68;
mem[16'hFDFD] = 8'hA4;
mem[16'hFDFE] = 8'h35;
mem[16'hFDFF] = 8'h60;
mem[16'hFE00] = 8'hC6;
mem[16'hFE01] = 8'h34;
mem[16'hFE02] = 8'hF0;
mem[16'hFE03] = 8'h9F;
mem[16'hFE04] = 8'hCA;
mem[16'hFE05] = 8'hD0;
mem[16'hFE06] = 8'h16;
mem[16'hFE07] = 8'hC9;
mem[16'hFE08] = 8'hBA;
mem[16'hFE09] = 8'hD0;
mem[16'hFE0A] = 8'hBB;
mem[16'hFE0B] = 8'h85;
mem[16'hFE0C] = 8'h31;
mem[16'hFE0D] = 8'hA5;
mem[16'hFE0E] = 8'h3E;
mem[16'hFE0F] = 8'h91;
mem[16'hFE10] = 8'h40;
mem[16'hFE11] = 8'hE6;
mem[16'hFE12] = 8'h40;
mem[16'hFE13] = 8'hD0;
mem[16'hFE14] = 8'h02;
mem[16'hFE15] = 8'hE6;
mem[16'hFE16] = 8'h41;
mem[16'hFE17] = 8'h60;
mem[16'hFE18] = 8'hA4;
mem[16'hFE19] = 8'h34;
mem[16'hFE1A] = 8'hB9;
mem[16'hFE1B] = 8'hFF;
mem[16'hFE1C] = 8'h01;
mem[16'hFE1D] = 8'h85;
mem[16'hFE1E] = 8'h31;
mem[16'hFE1F] = 8'h60;
mem[16'hFE20] = 8'hA2;
mem[16'hFE21] = 8'h01;
mem[16'hFE22] = 8'hB5;
mem[16'hFE23] = 8'h3E;
mem[16'hFE24] = 8'h95;
mem[16'hFE25] = 8'h42;
mem[16'hFE26] = 8'h95;
mem[16'hFE27] = 8'h44;
mem[16'hFE28] = 8'hCA;
mem[16'hFE29] = 8'h10;
mem[16'hFE2A] = 8'hF7;
mem[16'hFE2B] = 8'h60;
mem[16'hFE2C] = 8'hB1;
mem[16'hFE2D] = 8'h3C;
mem[16'hFE2E] = 8'h91;
mem[16'hFE2F] = 8'h42;
mem[16'hFE30] = 8'h20;
mem[16'hFE31] = 8'hB4;
mem[16'hFE32] = 8'hFC;
mem[16'hFE33] = 8'h90;
mem[16'hFE34] = 8'hF7;
mem[16'hFE35] = 8'h60;
mem[16'hFE36] = 8'hB1;
mem[16'hFE37] = 8'h3C;
mem[16'hFE38] = 8'hD1;
mem[16'hFE39] = 8'h42;
mem[16'hFE3A] = 8'hF0;
mem[16'hFE3B] = 8'h1C;
mem[16'hFE3C] = 8'h20;
mem[16'hFE3D] = 8'h92;
mem[16'hFE3E] = 8'hFD;
mem[16'hFE3F] = 8'hB1;
mem[16'hFE40] = 8'h3C;
mem[16'hFE41] = 8'h20;
mem[16'hFE42] = 8'hDA;
mem[16'hFE43] = 8'hFD;
mem[16'hFE44] = 8'hA9;
mem[16'hFE45] = 8'hA0;
mem[16'hFE46] = 8'h20;
mem[16'hFE47] = 8'hED;
mem[16'hFE48] = 8'hFD;
mem[16'hFE49] = 8'hA9;
mem[16'hFE4A] = 8'hA8;
mem[16'hFE4B] = 8'h20;
mem[16'hFE4C] = 8'hED;
mem[16'hFE4D] = 8'hFD;
mem[16'hFE4E] = 8'hB1;
mem[16'hFE4F] = 8'h42;
mem[16'hFE50] = 8'h20;
mem[16'hFE51] = 8'hDA;
mem[16'hFE52] = 8'hFD;
mem[16'hFE53] = 8'hA9;
mem[16'hFE54] = 8'hA9;
mem[16'hFE55] = 8'h20;
mem[16'hFE56] = 8'hED;
mem[16'hFE57] = 8'hFD;
mem[16'hFE58] = 8'h20;
mem[16'hFE59] = 8'hB4;
mem[16'hFE5A] = 8'hFC;
mem[16'hFE5B] = 8'h90;
mem[16'hFE5C] = 8'hD9;
mem[16'hFE5D] = 8'h60;
mem[16'hFE5E] = 8'h20;
mem[16'hFE5F] = 8'h75;
mem[16'hFE60] = 8'hFE;
mem[16'hFE61] = 8'hA9;
mem[16'hFE62] = 8'h14;
mem[16'hFE63] = 8'h48;
mem[16'hFE64] = 8'h20;
mem[16'hFE65] = 8'hD0;
mem[16'hFE66] = 8'hF8;
mem[16'hFE67] = 8'h20;
mem[16'hFE68] = 8'h53;
mem[16'hFE69] = 8'hF9;
mem[16'hFE6A] = 8'h85;
mem[16'hFE6B] = 8'h3A;
mem[16'hFE6C] = 8'h84;
mem[16'hFE6D] = 8'h3B;
mem[16'hFE6E] = 8'h68;
mem[16'hFE6F] = 8'h38;
mem[16'hFE70] = 8'hE9;
mem[16'hFE71] = 8'h01;
mem[16'hFE72] = 8'hD0;
mem[16'hFE73] = 8'hEF;
mem[16'hFE74] = 8'h60;
mem[16'hFE75] = 8'h8A;
mem[16'hFE76] = 8'hF0;
mem[16'hFE77] = 8'h07;
mem[16'hFE78] = 8'hB5;
mem[16'hFE79] = 8'h3C;
mem[16'hFE7A] = 8'h95;
mem[16'hFE7B] = 8'h3A;
mem[16'hFE7C] = 8'hCA;
mem[16'hFE7D] = 8'h10;
mem[16'hFE7E] = 8'hF9;
mem[16'hFE7F] = 8'h60;
mem[16'hFE80] = 8'hA0;
mem[16'hFE81] = 8'h3F;
mem[16'hFE82] = 8'hD0;
mem[16'hFE83] = 8'h02;
mem[16'hFE84] = 8'hA0;
mem[16'hFE85] = 8'hFF;
mem[16'hFE86] = 8'h84;
mem[16'hFE87] = 8'h32;
mem[16'hFE88] = 8'h60;
mem[16'hFE89] = 8'hA9;
mem[16'hFE8A] = 8'h00;
mem[16'hFE8B] = 8'h85;
mem[16'hFE8C] = 8'h3E;
mem[16'hFE8D] = 8'hA2;
mem[16'hFE8E] = 8'h38;
mem[16'hFE8F] = 8'hA0;
mem[16'hFE90] = 8'h1B;
mem[16'hFE91] = 8'hD0;
mem[16'hFE92] = 8'h08;
mem[16'hFE93] = 8'hA9;
mem[16'hFE94] = 8'h00;
mem[16'hFE95] = 8'h85;
mem[16'hFE96] = 8'h3E;
mem[16'hFE97] = 8'hA2;
mem[16'hFE98] = 8'h36;
mem[16'hFE99] = 8'hA0;
mem[16'hFE9A] = 8'hF0;
mem[16'hFE9B] = 8'hA5;
mem[16'hFE9C] = 8'h3E;
mem[16'hFE9D] = 8'h29;
mem[16'hFE9E] = 8'h0F;
mem[16'hFE9F] = 8'hF0;
mem[16'hFEA0] = 8'h06;
mem[16'hFEA1] = 8'h09;
mem[16'hFEA2] = 8'hC0;
mem[16'hFEA3] = 8'hA0;
mem[16'hFEA4] = 8'h00;
mem[16'hFEA5] = 8'hF0;
mem[16'hFEA6] = 8'h02;
mem[16'hFEA7] = 8'hA9;
mem[16'hFEA8] = 8'hFD;
mem[16'hFEA9] = 8'h94;
mem[16'hFEAA] = 8'h00;
mem[16'hFEAB] = 8'h95;
mem[16'hFEAC] = 8'h01;
mem[16'hFEAD] = 8'h60;
mem[16'hFEAE] = 8'hEA;
mem[16'hFEAF] = 8'hD1;
mem[16'hFEB0] = 8'h4C;
mem[16'hFEB1] = 8'h00;
mem[16'hFEB2] = 8'hE0;
mem[16'hFEB3] = 8'h4C;
mem[16'hFEB4] = 8'h03;
mem[16'hFEB5] = 8'hE0;
mem[16'hFEB6] = 8'h20;
mem[16'hFEB7] = 8'h75;
mem[16'hFEB8] = 8'hFE;
mem[16'hFEB9] = 8'h20;
mem[16'hFEBA] = 8'h3F;
mem[16'hFEBB] = 8'hFF;
mem[16'hFEBC] = 8'h6C;
mem[16'hFEBD] = 8'h3A;
mem[16'hFEBE] = 8'h00;
mem[16'hFEBF] = 8'h4C;
mem[16'hFEC0] = 8'hD7;
mem[16'hFEC1] = 8'hFA;
mem[16'hFEC2] = 8'h60;
mem[16'hFEC3] = 8'hEA;
mem[16'hFEC4] = 8'h60;
mem[16'hFEC5] = 8'hC2;
mem[16'hFEC6] = 8'hF2;
mem[16'hFEC7] = 8'hF9;
mem[16'hFEC8] = 8'hE1;
mem[16'hFEC9] = 8'hEE;
mem[16'hFECA] = 8'h4C;
mem[16'hFECB] = 8'hF8;
mem[16'hFECC] = 8'h03;
mem[16'hFECD] = 8'hA9;
mem[16'hFECE] = 8'h40;
mem[16'hFECF] = 8'h20;
mem[16'hFED0] = 8'hC9;
mem[16'hFED1] = 8'hFC;
mem[16'hFED2] = 8'hA0;
mem[16'hFED3] = 8'h27;
mem[16'hFED4] = 8'hA2;
mem[16'hFED5] = 8'h00;
mem[16'hFED6] = 8'h41;
mem[16'hFED7] = 8'h3C;
mem[16'hFED8] = 8'h48;
mem[16'hFED9] = 8'hA1;
mem[16'hFEDA] = 8'h3C;
mem[16'hFEDB] = 8'h20;
mem[16'hFEDC] = 8'hED;
mem[16'hFEDD] = 8'hFE;
mem[16'hFEDE] = 8'h20;
mem[16'hFEDF] = 8'hBA;
mem[16'hFEE0] = 8'hFC;
mem[16'hFEE1] = 8'hA0;
mem[16'hFEE2] = 8'h1D;
mem[16'hFEE3] = 8'h68;
mem[16'hFEE4] = 8'h90;
mem[16'hFEE5] = 8'hEE;
mem[16'hFEE6] = 8'hA0;
mem[16'hFEE7] = 8'h22;
mem[16'hFEE8] = 8'h20;
mem[16'hFEE9] = 8'hED;
mem[16'hFEEA] = 8'hFE;
mem[16'hFEEB] = 8'hF0;
mem[16'hFEEC] = 8'h4D;
mem[16'hFEED] = 8'hA2;
mem[16'hFEEE] = 8'h10;
mem[16'hFEEF] = 8'h0A;
mem[16'hFEF0] = 8'h20;
mem[16'hFEF1] = 8'hD6;
mem[16'hFEF2] = 8'hFC;
mem[16'hFEF3] = 8'hD0;
mem[16'hFEF4] = 8'hFA;
mem[16'hFEF5] = 8'h60;
mem[16'hFEF6] = 8'h20;
mem[16'hFEF7] = 8'h00;
mem[16'hFEF8] = 8'hFE;
mem[16'hFEF9] = 8'h68;
mem[16'hFEFA] = 8'h68;
mem[16'hFEFB] = 8'hD0;
mem[16'hFEFC] = 8'h6C;
mem[16'hFEFD] = 8'h20;
mem[16'hFEFE] = 8'hFA;
mem[16'hFEFF] = 8'hFC;
mem[16'hFF00] = 8'hA9;
mem[16'hFF01] = 8'h16;
mem[16'hFF02] = 8'h20;
mem[16'hFF03] = 8'hC9;
mem[16'hFF04] = 8'hFC;
mem[16'hFF05] = 8'h85;
mem[16'hFF06] = 8'h2E;
mem[16'hFF07] = 8'h20;
mem[16'hFF08] = 8'hFA;
mem[16'hFF09] = 8'hFC;
mem[16'hFF0A] = 8'hA0;
mem[16'hFF0B] = 8'h24;
mem[16'hFF0C] = 8'h20;
mem[16'hFF0D] = 8'hFD;
mem[16'hFF0E] = 8'hFC;
mem[16'hFF0F] = 8'hB0;
mem[16'hFF10] = 8'hF9;
mem[16'hFF11] = 8'h20;
mem[16'hFF12] = 8'hFD;
mem[16'hFF13] = 8'hFC;
mem[16'hFF14] = 8'hA0;
mem[16'hFF15] = 8'h3B;
mem[16'hFF16] = 8'h20;
mem[16'hFF17] = 8'hEC;
mem[16'hFF18] = 8'hFC;
mem[16'hFF19] = 8'h81;
mem[16'hFF1A] = 8'h3C;
mem[16'hFF1B] = 8'h45;
mem[16'hFF1C] = 8'h2E;
mem[16'hFF1D] = 8'h85;
mem[16'hFF1E] = 8'h2E;
mem[16'hFF1F] = 8'h20;
mem[16'hFF20] = 8'hBA;
mem[16'hFF21] = 8'hFC;
mem[16'hFF22] = 8'hA0;
mem[16'hFF23] = 8'h35;
mem[16'hFF24] = 8'h90;
mem[16'hFF25] = 8'hF0;
mem[16'hFF26] = 8'h20;
mem[16'hFF27] = 8'hEC;
mem[16'hFF28] = 8'hFC;
mem[16'hFF29] = 8'hC5;
mem[16'hFF2A] = 8'h2E;
mem[16'hFF2B] = 8'hF0;
mem[16'hFF2C] = 8'h0D;
mem[16'hFF2D] = 8'hA9;
mem[16'hFF2E] = 8'hC5;
mem[16'hFF2F] = 8'h20;
mem[16'hFF30] = 8'hED;
mem[16'hFF31] = 8'hFD;
mem[16'hFF32] = 8'hA9;
mem[16'hFF33] = 8'hD2;
mem[16'hFF34] = 8'h20;
mem[16'hFF35] = 8'hED;
mem[16'hFF36] = 8'hFD;
mem[16'hFF37] = 8'h20;
mem[16'hFF38] = 8'hED;
mem[16'hFF39] = 8'hFD;
mem[16'hFF3A] = 8'hA9;
mem[16'hFF3B] = 8'h87;
mem[16'hFF3C] = 8'h4C;
mem[16'hFF3D] = 8'hED;
mem[16'hFF3E] = 8'hFD;
mem[16'hFF3F] = 8'hA5;
mem[16'hFF40] = 8'h48;
mem[16'hFF41] = 8'h48;
mem[16'hFF42] = 8'hA5;
mem[16'hFF43] = 8'h45;
mem[16'hFF44] = 8'hA6;
mem[16'hFF45] = 8'h46;
mem[16'hFF46] = 8'hA4;
mem[16'hFF47] = 8'h47;
mem[16'hFF48] = 8'h28;
mem[16'hFF49] = 8'h60;
mem[16'hFF4A] = 8'h85;
mem[16'hFF4B] = 8'h45;
mem[16'hFF4C] = 8'h86;
mem[16'hFF4D] = 8'h46;
mem[16'hFF4E] = 8'h84;
mem[16'hFF4F] = 8'h47;
mem[16'hFF50] = 8'h08;
mem[16'hFF51] = 8'h68;
mem[16'hFF52] = 8'h85;
mem[16'hFF53] = 8'h48;
mem[16'hFF54] = 8'hBA;
mem[16'hFF55] = 8'h86;
mem[16'hFF56] = 8'h49;
mem[16'hFF57] = 8'hD8;
mem[16'hFF58] = 8'h60;
mem[16'hFF59] = 8'h20;
mem[16'hFF5A] = 8'h84;
mem[16'hFF5B] = 8'hFE;
mem[16'hFF5C] = 8'h20;
mem[16'hFF5D] = 8'h2F;
mem[16'hFF5E] = 8'hFB;
mem[16'hFF5F] = 8'h20;
mem[16'hFF60] = 8'h93;
mem[16'hFF61] = 8'hFE;
mem[16'hFF62] = 8'h20;
mem[16'hFF63] = 8'h89;
mem[16'hFF64] = 8'hFE;
mem[16'hFF65] = 8'hD8;
mem[16'hFF66] = 8'h20;
mem[16'hFF67] = 8'h3A;
mem[16'hFF68] = 8'hFF;
mem[16'hFF69] = 8'hA9;
mem[16'hFF6A] = 8'hAA;
mem[16'hFF6B] = 8'h85;
mem[16'hFF6C] = 8'h33;
mem[16'hFF6D] = 8'h20;
mem[16'hFF6E] = 8'h67;
mem[16'hFF6F] = 8'hFD;
mem[16'hFF70] = 8'h20;
mem[16'hFF71] = 8'hC7;
mem[16'hFF72] = 8'hFF;
mem[16'hFF73] = 8'h20;
mem[16'hFF74] = 8'hA7;
mem[16'hFF75] = 8'hFF;
mem[16'hFF76] = 8'h84;
mem[16'hFF77] = 8'h34;
mem[16'hFF78] = 8'hA0;
mem[16'hFF79] = 8'h17;
mem[16'hFF7A] = 8'h88;
mem[16'hFF7B] = 8'h30;
mem[16'hFF7C] = 8'hE8;
mem[16'hFF7D] = 8'hD9;
mem[16'hFF7E] = 8'hCC;
mem[16'hFF7F] = 8'hFF;
mem[16'hFF80] = 8'hD0;
mem[16'hFF81] = 8'hF8;
mem[16'hFF82] = 8'h20;
mem[16'hFF83] = 8'hBE;
mem[16'hFF84] = 8'hFF;
mem[16'hFF85] = 8'hA4;
mem[16'hFF86] = 8'h34;
mem[16'hFF87] = 8'h4C;
mem[16'hFF88] = 8'h73;
mem[16'hFF89] = 8'hFF;
mem[16'hFF8A] = 8'hA2;
mem[16'hFF8B] = 8'h03;
mem[16'hFF8C] = 8'h0A;
mem[16'hFF8D] = 8'h0A;
mem[16'hFF8E] = 8'h0A;
mem[16'hFF8F] = 8'h0A;
mem[16'hFF90] = 8'h0A;
mem[16'hFF91] = 8'h26;
mem[16'hFF92] = 8'h3E;
mem[16'hFF93] = 8'h26;
mem[16'hFF94] = 8'h3F;
mem[16'hFF95] = 8'hCA;
mem[16'hFF96] = 8'h10;
mem[16'hFF97] = 8'hF8;
mem[16'hFF98] = 8'hA5;
mem[16'hFF99] = 8'h31;
mem[16'hFF9A] = 8'hD0;
mem[16'hFF9B] = 8'h06;
mem[16'hFF9C] = 8'hB5;
mem[16'hFF9D] = 8'h3F;
mem[16'hFF9E] = 8'h95;
mem[16'hFF9F] = 8'h3D;
mem[16'hFFA0] = 8'h95;
mem[16'hFFA1] = 8'h41;
mem[16'hFFA2] = 8'hE8;
mem[16'hFFA3] = 8'hF0;
mem[16'hFFA4] = 8'hF3;
mem[16'hFFA5] = 8'hD0;
mem[16'hFFA6] = 8'h06;
mem[16'hFFA7] = 8'hA2;
mem[16'hFFA8] = 8'h00;
mem[16'hFFA9] = 8'h86;
mem[16'hFFAA] = 8'h3E;
mem[16'hFFAB] = 8'h86;
mem[16'hFFAC] = 8'h3F;
mem[16'hFFAD] = 8'hB9;
mem[16'hFFAE] = 8'h00;
mem[16'hFFAF] = 8'h02;
mem[16'hFFB0] = 8'hC8;
mem[16'hFFB1] = 8'h49;
mem[16'hFFB2] = 8'hB0;
mem[16'hFFB3] = 8'hC9;
mem[16'hFFB4] = 8'h0A;
mem[16'hFFB5] = 8'h90;
mem[16'hFFB6] = 8'hD3;
mem[16'hFFB7] = 8'h69;
mem[16'hFFB8] = 8'h88;
mem[16'hFFB9] = 8'hC9;
mem[16'hFFBA] = 8'hFA;
mem[16'hFFBB] = 8'hB0;
mem[16'hFFBC] = 8'hCD;
mem[16'hFFBD] = 8'h60;
mem[16'hFFBE] = 8'hA9;
mem[16'hFFBF] = 8'hFE;
mem[16'hFFC0] = 8'h48;
mem[16'hFFC1] = 8'hB9;
mem[16'hFFC2] = 8'hE3;
mem[16'hFFC3] = 8'hFF;
mem[16'hFFC4] = 8'h48;
mem[16'hFFC5] = 8'hA5;
mem[16'hFFC6] = 8'h31;
mem[16'hFFC7] = 8'hA0;
mem[16'hFFC8] = 8'h00;
mem[16'hFFC9] = 8'h84;
mem[16'hFFCA] = 8'h31;
mem[16'hFFCB] = 8'h60;
mem[16'hFFCC] = 8'hBC;
mem[16'hFFCD] = 8'hB2;
mem[16'hFFCE] = 8'hBE;
mem[16'hFFCF] = 8'hB2;
mem[16'hFFD0] = 8'hEF;
mem[16'hFFD1] = 8'hC4;
mem[16'hFFD2] = 8'hB2;
mem[16'hFFD3] = 8'hA9;
mem[16'hFFD4] = 8'hBB;
mem[16'hFFD5] = 8'hA6;
mem[16'hFFD6] = 8'hA4;
mem[16'hFFD7] = 8'h06;
mem[16'hFFD8] = 8'h95;
mem[16'hFFD9] = 8'h07;
mem[16'hFFDA] = 8'h02;
mem[16'hFFDB] = 8'h05;
mem[16'hFFDC] = 8'hF0;
mem[16'hFFDD] = 8'h00;
mem[16'hFFDE] = 8'hEB;
mem[16'hFFDF] = 8'h93;
mem[16'hFFE0] = 8'hA7;
mem[16'hFFE1] = 8'hC6;
mem[16'hFFE2] = 8'h99;
mem[16'hFFE3] = 8'hB2;
mem[16'hFFE4] = 8'hC9;
mem[16'hFFE5] = 8'hBE;
mem[16'hFFE6] = 8'hC1;
mem[16'hFFE7] = 8'h35;
mem[16'hFFE8] = 8'h8C;
mem[16'hFFE9] = 8'hC4;
mem[16'hFFEA] = 8'h96;
mem[16'hFFEB] = 8'hAF;
mem[16'hFFEC] = 8'h17;
mem[16'hFFED] = 8'h17;
mem[16'hFFEE] = 8'h2B;
mem[16'hFFEF] = 8'h1F;
mem[16'hFFF0] = 8'h83;
mem[16'hFFF1] = 8'h7F;
mem[16'hFFF2] = 8'h5D;
mem[16'hFFF3] = 8'hCC;
mem[16'hFFF4] = 8'hB5;
mem[16'hFFF5] = 8'hFC;
mem[16'hFFF6] = 8'h17;
mem[16'hFFF7] = 8'h17;
mem[16'hFFF8] = 8'hF5;
mem[16'hFFF9] = 8'h03;
mem[16'hFFFA] = 8'hFB;
mem[16'hFFFB] = 8'h03;
mem[16'hFFFC] = 8'hB6;
mem[16'hFFFD] = 8'h8E;
mem[16'hFFFE] = 8'h40;
mem[16'hFFFF] = 8'hFA;
  end

endmodule